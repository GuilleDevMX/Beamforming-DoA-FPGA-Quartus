��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���~�`���sB�U	Ù���iCK�������Kuy�y�	���5r~��O*�7+�[�r�E����Y���5K��y|_,�A���d�+!�c�����mk�_v�c�O;F�@��3�s*b��	�O|r��d�gG��-�
�y�Nh��4G���Z�;x�����S�I��r�����1	��L&��I��%
;td\,��_�I�)��������]�x�9�u�Y0U�A�EB�B��.E����Ƽ�Y�F>h�f���8��g��� J~MJ�l��Kt�>��-^x��<�\�sn =e�[#Jǭ�%^O��e3g{y+&{f�c{��"CV�Y��+�M9��/�<��m�1q����L��̊�.�v�Ā)n2�2bO�!�����ǳT�6�z�0��TiX�]��c��[8�2/jn�9L^J'��gE��^;g���U�M$,"ʇETb�\U<'��eC�1�~]��H��2���T�]ہ��B���
}�m��'7m�!�l�f��W�:�L%�A�^��e�Y���>�nA"3�x4�^ lR|&䞈�An��q���Z]�ȉ�閇G��A	W��d&�r~��@ye9�4j��u��*o�C�_�>w��J�FׁAJ��p{&�
_��2�T�ϲn�gb���I��0>�3`�b?UH��yd���Z�|h��u�Pr���b����y�4W4ޥ3~��8:xt������:��Ô��<x��٫�z ����,�xG{o;`�p|�����I샪���/-��roJo��hs �����w�� ��Q;~ҝ
��{!	�v�I����s/\2�@&�Ol�O5Y�s��N�l!��t=)�s�N$��B�U��C#v�^�\���[nܷ/%X�L�ag? ���<��g�dY�:�&���kx��`O��l�,�]�o���
̓O^�{Ä��f��;�M3DI�L�����P:�\�?e/Oڱ����b4���gr�7�3Oz�:v
���\�W�K�.��f�P����/�	�1U˒6K P�����y��������~��L�&u�-	����ֹ�0AAFT��(��H���ֲױ~-��%���>��ӧc��T�/Tg R
��2;]a���"�i��"�a�H��\R�ܞ�O�I��Z�Ig��YC��]��	��ư��;�1]��S�j]~6���aW�"V��6�r��Q����B��u�L�"�X\Hw�o�HGl�c<����+Ì��f�F�|#_����DH7�0G @�U�Ītc�T�*�&&d/�3�~��PɎqLB�f�R
�vt�B�C����ꡖR0HBw �L�r��)�j��L��*�F�OO�Mi�?��Ѽ��ʴ
��_��j[>�Cf�i�ښ0̎���<�:���X=.��m7*Ơ<���0�(P��̊X�|�C�1(�}���m�J B2W��P�E �b��F--�Zk�"8�:�\g3`㿑?��5���4��A��'g|"@�	�[������]��^I�]s��I����['+֚�� :���;�J�[�'�\H���1��Lϳ�\�R�+���*V�+��]��zV������Hb#-���.��O�������:[�>$�i��-ay_2�o-~������q^z�W��Ӷ���+��e�9^��p�͝:4(���q��D8S�]�c�/D����cT���>�ː�M��QUq�l(�By7��1(��-死��hL�	�kK�b��)-P.���*��f�]y�m��� V��,��� �5qM}�LK�V�\�a=��N �U��s<٣���<����l���[����%O�G�����+1(��o�_���:���{t�:Ί�ič��V�t*Yy�u�����q�g8:a�:é�`����Ά���O)0p�*�S��J;�5i��o�x�r`�J7�ׯ6<P�C�SR��>	�%I��|��ґP�6���M��c^I!��:3��f\A����m�S�쪑ý�6�,��k��$S�2�H��܇�~U>,98-k��R0S�-�