��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#u�.!�N����Y��%��ۈy���BV� �e�_�LTP�m1j�\��s�/ٝi[����H��'��x0Մ����H<l8��'ƹ��{�,u���x��%.P�Ʒ��;��צ�5��gt�3�/�O!)�����4��һ� ��{�s֨�}#�b��у�m?N<9x�9�a��1h%��S� G`���ao~��c5m�n�h�J+�rt�4e����l�d3I��[��G�:�N�;��б3��Rf&jS�ʼ3��<�zDM�7�ɢ����&�S�~�����;QY�ý���X����;�B���.��tȾ��ic��8/G?�^�>f�U���"��:=������`�J�1�71/��a�)lH�J��r~�:��I��i�cK���ѷ�[i��� �MndF�׻�3��$y��%lp9�� �m {�ş�`T&v�6.q���*:��r`�lm*��}�rl`��Y;:D��ش�Ń$��=�ނ�>5�|?ZtM�hC5�M��V"���jj`?��2h~�m-{f��e��l,�kLZ�tMf����k`�=P��B p(�]z*��c��� ��#0K��7f[~Tȴ��^���z��t�q���M��cw��9����n=%� �����������O$w}i�Nz>9v�C4�`Ӆ!$:�Aؼ��Y��j�S�z�q�H݃0�fl�	���B�yA8+l��;+���/;���S�S�#��$�Ө��Ȏ{ldluR�ם/`>%�7��(�3��������� �6�ު���;5ۉ\{��-�=�����%�飡gJ�� �PI�`�4���xߩ�B�7���2�C��΁��r���,��ݧ��]�8N� �	��'.��"�^�#��w!h��D��>����p�SҊ�G�)�5���TS�����eu@����T
��,�s;����j`����G®m��������TW�S�5Y�r&7l����z�xTh0��Ŗ�	�.��=#VqDO���@��@j�1=�6K)<V���`�*z~A��բ���XPr�ɘӐ=�0C�w�!��#r��r� !+�[�\5�Չ'�@��{9C��7�FƇ��g�an*'�w�-��k�� ���-�XeE�rI~���|�e�햒S�8������_T�^_}�bQQ�Ӻ��L��������]��"Z� �-�7o(҆�wlJ����S:�w����^�J�6�Eɮ���8���B0P˽�����}�Ut�ՒUvԙ�x)�}�*�_	rΘ%�F����.��W����4�k����f-�f�(�:�1�}Q!S���	�|F��`S����=fz����<S��qަ�^�Vf�n���~+O�F%����0n��Mm+�G�V%@�˹�z�����߷�=��l5@2�����Olb-���w�2��-5)����C��:CW��X3o��X��υ�Oͳ�I�9��W����L�/�I�'p��D��Aq^�Z�� �!ǐ������2A��\��@��	FcW8L&{��I��a�x7��FL���|w���qj����?����V��lJ(V賓�u3��༗Aq\k�>�� �s�^s��%�fp��8���������9<	jL�/h⓵�Z
����t�^L2���v��aq�g+u䀻�$Ll,���fKX�+�;�}F���)4������+9����
:.`� �[��ދ��W��En�	IـWtN)\�����#�����1��+�#�F>��i!\T�_S�F�������B�b��`3}�P0�/'ɗD��a����1�x��!���6䜮L��V���[���t�ر��]];	@!jT?������_��Q���l�9�^�$.�$uq��^ �0��y)k�3�S�"���2���4�a�P�o��B�0Y$����`/�b'˿Bρ�]M�������Ch1����"����`��ö���8���+Tyy��ah%tz�KJ���pp<�G��Y2�jkƏ�`�����R�ٌ�ES\nL%!1'Ź8_�x�0U��"�n\=�A=0�g#H�}�w�h�P*D�i�p�L��X\�;��n>~�F��R.�e24�9'�b���*ѽ=�+�gײ�j$ $=ox����z��T%' ��W�x�����U�yo����"��|�Qm��{c�;w�y���g{+�;~2 <)�_P�I��qu����:�JFgC�s-�-��]�s�e�����!�:���~���{�������59�����̏����q%r�ʰ�N��g0eދ�t��-�R��qR��b� ����͆T���n�5�7��Z��K�6� [��W*|��̓j0����%S�g%^)خ|ɕ����J���Q��@`�R���eY�~�XT�h�[fr�m��û������L42�Gc�����8����i�F���D��3��ʓ��h72�ֽݬ�Ś<�E�����kh�Q+���|�fJ�>�4QPv��}����,�V�/E�V�B���.�;&�.�=��Ó[#]�v� ��n�p
򁒾�ի`��RӀN��m����T��(x�k�<��	�f����X%���۾X�I!��"���)�<��� T���VM�b��>�YJ�1LL�_	j��:�eS�^eFvʴ�>'R�?�k`�(PF���8��I����S���F��#m�OŻ*��k"�)�mn��
@��ڀI�FK�3���d�Lۼ4��;ĭ�m��m�P��T.{t��"OOX#p���/fS�M�vJ�Ni�����/P\<��N�ƒU:���AX��s�QO@>��@�c�Զҥ�|�1XCE����V�:J���T�\N��M��7��?}ϐ�aƼ+=�~r��s��wmY@�C�x�}»����<�3��q%�)�Rp?�G��>�VA{�h�n��e�]���&ﯙ�*�I�OĞ��Fb�y0�$*<77�S9�M��\�� �m�v��)�%�I9�!	� ���P93<s\� �!YQ���2�f9/�uiA��m2 ��@��|��o�]k�99�?�Pᚽ���O��Z&�0��ۄ�RΣ�/V��l7������Jwr�D7.=�I�_��va_
�Ă���H�`7û~\d�$p$�~:��i��r�[�}�?��b�\����I�hI�CA�p��-B��������cx2x�xEC��o.}���렲^�߷��+���0�|�Xup��*5�	f+Uĝ�!�jע����	�6��p��ؓ��G8��*4�e�m���<@�p�>�x�Vr�	qF�ѧEY��x�7q�%�v�dh�����@i�i�I��3�4ݻ�ךZ^�)��٤M������Ge!Ň��o�:�|�
W��\��\�mIh��c�-�9��k��V����Wd��1�öGO.����.Q�u�_�K�Vv��q�oH.�N���mt͔��l�GwJ�����K��ZM����x���D�r@�_�����q�E~���jw�d��D+b�H�Ƈz�  g�\�}�4n YhD�����&9��r��zY��<̙��m�^�l�U�1�|d�.� �h�.F�N�]��7P���D_��0qa�!KR[�{_=�FpW�$8�._��f��N�YnVԶc0`Y��� �=��gh����U�)9m�0P���F���_^���3�2����*e���┹	�V�߱�L�s�BU�q��X���+��X���d8u�������LG[��1�`���V���%�J��<Ͼ�+02���ќ�]� ��?��x9�f�m-}&mx5�.?k���@��(����)S]8���ۊ%C����[��dM <Ֆ�=�f�l��U�[#e�ؿM�f��=�nK��=�2���E�:'���������!+�¢D�5[dMǕ��le��67 }f{�iֺ{���'����bd_�y��Fh��9���l�5Ua\t�!�'3�e�e�}�U�4]��.���9Y��رCHy[���b�2O��d�/���f����J��Yؠ~Uo�D6B�[��#��e)�]�녒�5��%d#0�#D����^�<a ��j�b9��%96�p@�I�Y�D���#95����g-(4Q���8i*���V?ȴ���u�����y�â�����&��9%V k?l�Kf��Gv~Y/�.,��9�Y��&ɼ[��G���[#� f"ܥE^)T٬��ayn����7sRw~%����H��;�Ð�^����( B8�R��A:�/T��K<�"��a�S$���ǘ^u���Ѝ�f� � XTX�1"�[�
�R˩����;�w1�02�d��?�+a�jga�pT.8���o����ym��T=7��[_5��O����_K#v��p�{�4<i�K�*/�Ft���4�-4��<�p����5[������g僡���<krW��P�p��<'�hwH@�r`�'��� ^��h�,�e/P³�c�GF�3�H��N&�'�[	�T�Ɏ��%&��w����	�{d�V���цaa��[-�906jk��"�>tޛ��Ɵ�<MJ�M˶�s/1�!>����s��8���C)V��	a�q�Տ��p�@�UWq0��5�0O�Z�T"BL��al�ٗz�)߾;��j��e y	����D�Zl{g	��+��ANxM�==��
Y�u�Ǯ�M�ˈ_����`�-��/%�<�{�=�WW��:&�`|�8;V*2G	ہ�;����08�o]bm��B��6>���*�"��"�DK�Ϡ��<H��&=�i��w�[D��l�}�:n�+�c�#��o�� m��@6��I�Y��"\u2*��O���/3�����Y�KVO�E�_co�o�2V"X-h+#�ׯ�!��u�h�em>*�8�@|�r�����>%o�0&���<��,��඗�mL�uGN��Ѯi�9����q����r���G�[/�eC�ZP��O#���	��Y���)L.\�Y����0꯲�Oe���w~jcQ��ԓ:���K��ϰ#�<��-�8x��)p������?�80�۠����c��6�m�_= H����i {����6n}$����<�B�����fOy�<bZ��
��'�#��X8�����[O��	���x+�W�.q>�%-ɼ�A�#���vJ|��kE��}�����`)�3���E&����w��I�O#<c̿#��r�^��W��k�-�O��;���<E66�d��ϳxN�q1�E�����(FR|����&6͵��?۴����\�j K��~5�7y�(LX:��z��óh���CBu�l�|�h.I��|���Ƨ�|A�B��I}Ϲ�ǎq���/� ��|>�������?y
�|�t�hB��B,�d�T��_`u�x��,3[dH�
U=X�A�@��N��0߫'hsg�������n�
��k��L��V���p�f��J[ �&uաѮ�Iބ�>�$z��Sy?��	��F	 �&��Z����VD���n�'Y�}����������W��J��N������8b�����<b��3|L�v���}ɨ�a�Wg%�s;�8r/�A6��ɺ�k�%�Й�q���,5�2��N��_Ʉ�Y�����?����Gܛ!�O�1�l
����7П�T96����*U��2�Ut]ڡ�m�����⫠E7�r(�/��|�;���.�଻���j�{������?lh����ʛ,�`N�lmy����{�@>D�v��P簡�|�N����{x��d��z�>��=u����������
;<�l�4��Ѷ�C���r���I�o9.���p}��)��Rce�j��B�s�\�E3z�G2�zK0c��Qo*�d)�=
�ڤ\����F?�@��m���&�W��F�.d�G-�q6Kr���
�����S�|��.�	m�!����u�R��)��.Z������d׍��<�X�)썔����w+��ހ�'��I!tM��MG��E���ɒf�a�i"��[�ɺ$��NP��yeM�e�W�82UŽ���}8�f�_	^F{&��#��l��n�G70�Ȃ���#� ���#�Wo�9\��1�ڧӬ��Vq�ӎ�L�V��؄�M��/s}�d\�?9�����%�P�)
E'�j�>�I&H�/E�E�+������'�2���nF&^>?���3}�8Fk
U ̕q��ے4�,�U`
I'��e����T�>�S�Ry�"�B�,FgfZ�ˀpF�f��;��h�L!����i��
ԺrNиF����NF�{���#?�a�7�����4!t��^i���,��q��2�7lzU�a[�w�$�oxv�*h�J���V��9���V�;;Ҫ5(��CO�i�6Z�Qp٧��QJXUYlc�e6s1<^&���[ˑ&�.>�=ψ�o��]��?�ʉ�K�%C����Y���� M��I�Xз#�bP�!iԜ�u���)n��i���� Y�D�ZIة�D
X��eu��_H��ʈ����r*Љ�./	0�+e� ����o�9x>���OI$$궁�
w@� ��v�_�C�����3��	�Q��y��"��"T�A�՜`��v�~�"]