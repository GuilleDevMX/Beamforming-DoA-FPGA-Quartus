��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C��(b�g L(� �?�ڸ���b?p~�����1��/5������'�#�R@~b^-d!,blCHa
���&'sDH���r�iJп��J��&��׎�GH�t��LP��7-o\�㱄~C6���k̜4�����m`��:���>>=��IU�	�Tv�e���)"���wӿ���u+=�Ux%��(��_�j�I^ƭ����'�*�ob>+�(ud��^�\kr}����I7��,��A�����9n{B�*x�"(��e�Ÿ�O�e]n�+�X��}�T*=�<�Tr�?@�N�j��H�[ڦb���a�%�ߛW��t�!º�^��j�u{��!VQ�)��{��k�Q,o]��n�'�qAZ�]��ȧ�Bgg0|[8��zJT�O$�vV�6��ʠ�w1Z�d�P}�d��Lr���)��0e�[��m�&Ԯm(`���T�a��.~=;��]��VM.=�Ni0DyJ�V���{�?8m�>e�'�]�+�E��L+��z=g�' ��ҐO'����:�Nxas}w�cs\G���;G!�?Ve!�����m�q|V�F.T�E��pTW�9��x�����nu�+����N���ZQ��h�,a�������~��PJ�x�����`�zO��͖��#~����M��e��w-Æ�(L@��58�=�ׄ��^�����4��U]���¦����*�̮,�<*<��࠽7�F�B���)��4��5MOe���b#M&�)Ҽ}ZҬ!y�Vj4Ȕ^Lg�%���: �9�'�N�F�7��^x�I�����{oU�U�}V�C�u������n5����-1E_�7��)V����N��"�4��#9ߊ���5-YI ���{?���h��8���
�Vy��z�]p�*���-����6�Q��(��4�ll�l#����f��I�"е��@�2�@#�`[��쐗ժ��u�����h�m�{/>���c/N�����Gs�.�D4��������g�x&��]��5��f���bDY4�	���yu<��F�����m]}�/2h&���h���GC�^�W�C���<y:���:0���vJ��#�"���1%Ӆgxi��9l��H�F�а�����g;\�#V]��.���_���=iۿWp�`����<}&<�*g_�<�Q�M`�cJY���CU�xX�j՟f�jn�80��Y"�6�Ɍ~Y�������K��M["Ҷ�sKI$ٛ'����Y^G_n6^kc���יT8�]�����d�x�������Y��iu��ޝJ��~Æ��`�Ջ�$��PS�p��"3@?B&�&�)����2��:A�� p����6�h����^��])��n'�	��bu+���@�?��A��|(C�#��W���zH��?��I�@jc�Ed��mq��E�D���K�J�t��,l���t� 6�߬5!N���1�`E�̬�~1��w'g�ކ�;�fi�)�'n��E�2�=��%�K�q4«�ed�
�^�̦�d����:t�����%tA��t��$5q�r^m��JT��Ao"���A2��$у3F�V���kt{�ty1@��^���F1�U�� �!3���v�]��e������p�S߀P���H���*K�(>��,�Ճ�/����F^Uq!� i��R$&��/�;x^%�o��"mX �/����M�))f��_-FD�x�iS�W�tB|悍k/�m��8��g0��T��1;�*�g�<���Z�^X��1�>Ż+�FD���0��d� ��'�=�q���{�ј�C���ZSܒ�r��v��H+���mɾy�k��!�~�*|�s;/�_�f3*��n��Y��O� ?q���Jh	m�}ij�[W#5`�Ψ���>��)%�x�n��!#�#/x����㴫���U�T�AF+ƣ�j���sjg �v�z���G+fz��m"�"�z��n�v�z��Ht�E����Dݳ�ލ2ٔ���d2]�uHjҀ!�aa���q=9ꙁϥ�;�=0��@���K��q�<������A���Q�5��ߊF�GJ�����8=2��"�'�4�"����4(����^����-3������_�-�t�K��m��WB"�N:r�Ň-8���v:*����,q8&Gآ]�ݜ�	���c��U�'@��R`����h�B� C������<�Fk���n�#�CE/����s@y>��s9@ <mg�j&��J��*(Ѻ�ɹu�fZ�>e�9J�O����g����8K�u5d�������}
�E`8���Pp�
��NI[wR�A���=0��!V$�d�ș�(�3yw�۞O]a��� /Вy�h	UQ��<����@$��p�~P��M���hX��]<r	��R�	&��A7_�H���<jD���g���p�xQ|�r�L�	�!����U�ڙ�"�R�+9g���""q/3m���q��@�p���Jk�,Ӛ���cH�NM1H�'�í��|��K�xy0RQ;�>�����	�9�i�k������U��WKA��/�O�8\~K��cpS"M*��W�F3P�.�h&x�'^��W���U󒫞J�>,���qW}.{4���33N�:8g��P�^`��{����k���{c���MҥXG����i��]�ו�����.F��8�0�������'��w�a`�l��J'I���>�I�Zk�P�-�^US�iy�+B�����S�F:��B�>��8���a�/�#B"G�;���Л�r6�ҰD�$�/-�E��iH^:�s�Xi��D-kn鋅�O��+ĵ��P�S`�