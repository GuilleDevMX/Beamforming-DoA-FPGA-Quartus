��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V��������H[H�6.�{Sh~>�>��v����E$	���Y~P��jc�Ƴ�7Q�|P�Y�\�y��S^Ḳ�$kK�PF����M&��uA��`Ne��?�Ի��������ou�&Yh��d��"#�; q����8�'��O�	Rv%�(��f�gz?7D��:��%���xhr>���aCs߿�d�@�0n��,;0��ؠ�s&Dϕ'��T�X�R���'�V�S�YjZlJ��K�HP#��
5�����Ǹ����å�wJ�h.����SlECށ��p�upMT�S�6�?W	)�Q�i;������'�X�VӚણ��q'�{��"�x�J9��bWbR�:J�O����~C0��w��5�j`|+#�F�޳4	������/_�T���H����(��Zle�F,Yn�ܺG�_���
UL*�DF�N�ش��%=��<Y�-�� ��T�D^�h�V��wn������Ӎ�[������a��I�?�h� ���(v3�d�ݐr]� g�����9�y9�Ϙ�*&�E錒�'�Jt韅���Cs=R�M ���3%Ǧ��k(
�|�n}��7�2���0f��,��ܭ�O^�]�@����;R�]=��t��>�9�$�����u	3L�l�h���#yX����z+�c����f_���\w�5�+&��=�����s�Pc��;K�5ڶ�S����.yv���;n<����nܖ���Q?]�jc�N\I�t��0��?Y�<δ�)����i@��SA �����p
�s���X0�W�5B����0��ɸiE��`w��Xl����I=^ǳ��q��� �F��r��3�o7eB�T�� ]Le�-#�uX���K_M�.<s��e��W�� �l�1j��f�9g������հ����'Ζr�r��LN����IB1���9��E����ڢ��G-�!W0�(�!E����R,k�,��CƉ��s��E�����Gr;��������
a1�R��*�@�#D#�/���N��$��Þt~W�p?��>���c\w���D�(�h�F�B�ʋ����v�%^��d+��y0`7~V���x����9N��"/��r�{`�\L.J�ehlp�טgֈ�!W2��<��2�,�	}������{�9ۋ�m�p�����3���ZBs�v� �����0��m4�)��Ml�FnFz���ב��h���g(�o��l�m݇N�;6^D�fs�2h�L�~��Q��7��E�,О�c��̨�J��546+d&Ͼ��W'7�.�� ��Q�@A���&�����c���ˊ�X�m�
���q:'�	o�.�$E�2���pX�<:�%�8Aq@C-�V�X䤩�(��}�t�e���|�2Ł�z���r����P(T���P �� �������)�-"�Ϗ�~=�����g)�*Q%+U"Z4���`%0�x�ʩ"��J���a�>=Ey��UJ�����J[��N�w��==\ ��3��;ȕH2B�0����f�4}fa٫��S�uyR���\?T�^�YP~L����ˁ7���T����ԻPRS�oF�(f]/�3��c��!���oR���UN�ܜ|�����"���D��QY�0�'f�K����L�{��jK��Q[�&
�ߣ����Hc }��feb^O�4����ڢw(p��鰑���Ɔ�8�8)b�؃�S��op`��
qk|��P��a;J�����+�Ev����s�kd4�>�H�L�7��V��&�>ē^�Q�6}��H<�h�0�<2`���w'���.��03����V�˿�%�f g�oX�ƨ�X �8�j���*P:�o9�a}Q��Gm�FE�sV�iN�����^���)B�u�����Jߋ�
�r�� �\̿���(^i��'���+��ը@ң�f�n��F���%����s�����v�����5L�.a�P���hP�'*y�i�-I�'~X��}��>s|�>n����΢���6����U���y��[cߛ�X=���-ԗ�)�J9}D�w�A���s/��:���w�X�\G7y�q.pVӊ�㑧�*�r}��U����$A��rm]j���F�Jx�{x�ȍ��N�}#�T�*�ي�N�Xĺ�	�s=@�N�'u"�W]g��T�n�Y]�z�PT�F����ϛeJ���/�&TY׫�����	��(�^PP�M�N5}��ރ0,�����-�!W�F2����L2�f�0H��Vk�XVY`��?��<�Ep�0�ۄ�`i �և��;wJܑ��tE ��]���Y͘^��ڗ)Y�&�]�t�k�}
{��;y���NnT�м���a�`���y�O�������ȵX�4�^:;|�����_����pl/�gS�ז�ː�S|��������=�=�k|T{��@�QA߾|Ew����$3-��T�x&��Zed 3+\�i	re.ݼ���2�B紽��r/�xp6�[�x{����=L޺ÿ(���ב��DػD5�`]O��D@ɟiʺ�ż|����Xs�$��D��I�K%C�g�_O:xN���jY���y�cp�;�=+�ZO�i�n7%[�$�֍�m�3�S�0[�'�	9FM�s�4��v�-y��j4���A�u��h�,+�	g��*m$�:��ow}Q��7���t�݋3ч�� �q�"�V��A��&	��-J!KT9q�5����m�u�aʄ0��B;Ȑ��G�Ƃm�t��Aa/M�~������.��Ș3ip�c��8~'[v���>�FT�Ö�bPx$�U{<A@����͗��fU޴�G�%��пd1+9���.J�����:%gw�a@V��1����t�2!�V�G(�k�P꥟pf���~`Iʏy�0Ĕ�	���W��5��ö�)>�<�[PD��v�}���{p9v
6��Stx���S��64�׍.Q�qVQ(i)��=��r��hX��fa����pCω��xY6��'�RR���Ө�}�O�$����|	ri-�BJG�����ْ�l&�`��!'ݯ��}���♫�L����M<��ù�9!����YA�vC��6�Tv�� W�z��x�f��K�}�b��^�G�ϤO�ٻ�L�|��Rh�H]S�p��f%��:��O��<��w�#�6�0�}/�?4�\���b����dw/s�G���{�X8�?v���EQ�c�>_m�������AZO���/]�
9��)�Q����1
�b���l�=���"�|"� ����\�as��iF3K}�H�V`n8U���:c�z�G��l�ơ���~��Sݩ᪫E%}�sϺ��Zh_���鬟�Z��#�Ö��/̳���wR}I��W�����Eĸ��8ciʣ��6�I�e�#s;bfM�"���h�b�j�,��Ar*jh���2�ڱ�Q��_e���8"۷�uҫo�B8�&�U�u�1�6�
��R����;aZ��L�^�J���v�)�6��o�7`K���ka��:����|L�V+��������t1�Q�*T�L��*�$��TG�e�N��d���Au�OE�?�"II�hA�(6�"�c�
F�)c-Zn��F?��^J�HCJV"ԭG9I�����*)�:�</�q����,	�Fj�C&�^ʵ�eݹl��q�H��h|o���R7=��U"��#v.�;�7c���cq�o�ck��l�q0q��Mk"}���E2ۗB�����#uU��R�s|ڏ�7�S����%Gi��v��p4K��7<��W3r_��e���͖�A�ON�{�O�ٻ"�:�*ڇ�änJh�R3�t��#� Q+��<׵+*w?PB%�u.�s�k��K���5��L��*�u9��S�25?1��A1?�ʝp��Z���b�y{ �J
�{���"im�`O�$g�a�j)��o���v7"F�W�d��z���M�.��`+q�R���|���W����'N�-3��/�G(
�=���J������Cg��y8|��QZԍ"���3Y?w7t��L�-yD�|�	D��"��p�v�+-����oĿ�z|��!Ǩ}Nx&��Q	5���U�n�k���15��T�/�����2�z�{|o�6s��ZR��NXK/ʅ�\�' �sƤ������N����&���φ  ;���e,���ذ�����Iǿe�@�rLg�j�? \ϴF�d�t�oƻ�;g�DA�݅�yX��US�xl2