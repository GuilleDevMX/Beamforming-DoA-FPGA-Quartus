��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���V�h�x���m��7�E�!�����s`*	v� �}]�73�Ƿ�-��u�9?Թ��̠���#�����'�Z=-�5�A+]�F�Օ?VjPH�`ҟ! ���-��*B��m�76�eu��r[&[��"��T�~A�H1v7|cQ�A[��n�`b�p�p���H៨0Z8�ٓ{g��W���"ǪMJ��F��S>@��j���-ČU�u0�!y�W�RԦ
~���x�S�7a6	|���-�U�>N�3�ޢ�I�n[9��v=Bx�[t{+�~9F�<�-���+�V�c��t���4�E8(a�����e	Y�΁���#z��˦[]'Y���b�B�ҿ���3]bN��n�Fn
߈� ���s��X2�a�.-n�v�D�&&���$T������[�:��p���V�į6�0E��s�����s7��"����|�=8(2:]$��l�<X��`&2�����I3�@:*?��%���@,}QB_4L"��}���oJ���?L9�����c"�v8� s�������2�J)��"EU|��0�Id<�D��π�{��I|p��0^;�x?��#���	�ZZ��U,7���lRЄg?A&���1Hĵ;l��>N�8:�qH_�yP%a�{�S�w@ū�p*����=8;=�ow�)�c�G�9�/n���
k�4�w1�u$��#ڍ�1`�.̭4jf���y�F����9��é�Ё�k�`9y��ͧk��,9�>����ۏ���*�1>�s�����%L�n����]<+8�i�����k�7˥Ob�Ϝ���ؕ�(�yK׽7X�j6���q'������?-.h�
aF�7A3'�Z�o�Hu�����
;���\�	�)ё���4gƧ�E�}���{pF�{�ْ,$ۼ�'f��ƞ�yR�yGT/a=�Z���NK���5�����a�?^�1=�<_�|ڧ#g��/M���r����v�3\:��O"ϟ�k
�A���ŧ����5J��^@�� 5ڌ���,�),#��>A-�l�){��ER|���������BL��	�}�u-����-/̶d��� ���+�*�����pmw������Egq��� ��!N�K�:I^�sQ;�T[�����&�U�X�/��*D���V���
~�anR�+w[��8�~Z��m�!��AǮ�ai�r�&���)��4�;_�E�o 9�Ӯ��]�M�6�kgwE ���?�ޞ���'O������Eع��m�,`�t�ό%3{��E��x[r�h��4�lǂK��z�b$�6��.����:`�oL��T�q?@f�0�p|`���\��ٹ��h�S�x�k7�z�a�`z�C����=���[��Gև�t���ֵMG�+����q�1�������� D2K��D1m=��ٹ�E���/�������늯�#?� R|�0�@
��,I��~��`J�d(�5ILy�v�hKe�ɑ1��H�{��w�����:Q���4S��!s�����N��"�)��=�&����y�����Z��qB#We��̉���E|^���$Nh0qk_ڷ�He��l�Ĭ��R����u�fE~��_�L�� �j�� �\/�Wp�MO���2F#ONs��-@ c��n�Ј���7<��2�W3u/j&Wg@Z�']��Giʁ�����M�3ԃ��Y�g��0���S�W�A��[5�IN3���.�e�<jz%~��!�.H��]�z�淍�(Ӷcc�?��/K�͚�������� ��a�-QӖ�����1�;_�a�9j��'�[�h4Js���-\�M��4P�?o����'��7ݸB��zcgO���a%��'��##f|���b��2/yA<���nJAt2���q������n1NB)�2�y�="��U��>ͱ'�SZ�n�*���!�l:��{�M`&��y�$u���5��q�N1��cr�Cr0���Xv(�����r3�-]}t��Z�2�f��_���f�{{�9m�dm�Q�]��X�׌��O�F�����ɒ*"�5m����i���A�|���oq
����2 x�w�'��A��}�b衿���K��A�������׍�]":o�C#ͯ��A�x��2�3�Z�ޱ�������>S�_/��n��-��E��Ñ��yn'[���+s��$�>ʶΪOu�O%nb�>\���i�Q{�U�m����i�5��%�J�]4�ˋ���ma��6��uU`	`��E�O#$�4D����K�����}��EѡH��d�����Q-2&g�5o�8H�y�m�܇�������{T��T<��v^�Ы���3�9egY$Y�����T9T���7�5N����i�</+n����9�T��aLUi�iw�4�VZ��q���Ϲ[���\���N0���>�T��.Dỷv�2}n<��%�^�C=C���ss��u��|��+�;F0��&�Y�=S*�l��v��(6^��D7�w���`�p�ۙN�0�`��;p��H,E���TMG/�#�n����{�U2dє�Y��-����@�N.ca8�b�	����b+�c���J���o��x;�,��ʜ/v�(3�)�N9�ph�2a0�t�|�J�އv��hf��@���2������HN�"O�\����W?_֛���B�F�(��Ç�ߏ8�z�I�)����Ȳ��u��Cjo6a!�I醮]ܗ1�
��W�6b}Ќ�@��Gh2����W���	�\�C�`|�f}g�'�{�O������9ほm�"l��B�n���Ϩ���M�������)i��j�<��O�[������Z�F��+�~�q̈́G=�v�|o�I-��o��K��]�� �OCF�?nk$�	|�w��&���,D�Nz-��T��ZV�^0�z������X�g#/��7�i:S �oAJA��_g���⑂�f�W;B��il���۴�W�W��6����:
)���=�d|S�¢�tཱི����6���mu�,QIzy*<�a��C~�F֢c��ȱ��?HU$P����5X_l<��)�V���&�wˤ��[�����D8Ӕ~�픿r!ԡ���eȊ�q�A�r����V^�`�R��$纺��p�(U-����6�;�2�9���J���5J�à�s=1���S7�N��&G&��u����w> \"�%����K��^)8���>���܂̖�T������x%\�O��=�N�'���X��ۮ������v�ɯ\-��8�|�1�%6ҧq��f$ڢڳiF�߷UaMLg�7Im�F�M W�ؘ�"�J���l����ն1��-ڮ����� U�ZO<?M�9�"�7��/����:)�����	��⟼O���K�i蔤>C�އ#�D+�O�uM="��G$\-��k������iy��g�=Q��jb�a�����#�h�73�D�I&�je��U���Y.�h{C<�`����8O</�!�P�f���D3I�m��E��ѧ���+�w �\��#+���P.���m���fz$2�8!B��U�����M!��X���h�w�t�:H�k�M��2�֎UKG$��,����
�w�bi����T�go(����b,�;;���f���́â5��3�G,]�����)�&f�\����J��[;$���ES��`����!�W� ��<^���Tѽ?#sk�T���1�B-5+�9!�X���>c���H��Oc`����k	�  9����Y��#Q��|Jhn��1t֩�*~-ƍ�50���g�:�?�{�]a�l�>�6��;(zUyw~l>�}� (�E����P�Ӂ	�0m�}����	Tx�
P��ii�~�~D\��k�'�?��{"9g3��|�F�+�|����V��{]�3���������L�v�J�${��rd䵜���y�]/!�d*mт���&ߟ���q^&�J%|��nX�ě�+,�5����Ky:�v�Y��1�`D��ʓ�����F�#N���`'�� �jVp4�=�.n_���1 &g�&�c�6<x����2��|ns0z�^���&��xy)9�%�WP��_�:J�O9��yz�(:��3J�'��Ox�D�`Q�4tUa`����I�0��\�_��s��?������e��X�$����֗��ƨ��}?���Ȩŝ-yQ$"�:.�̇ə��'bpw��ϕF���u�>lDY�ω���6c��ͭ���Kؓ+��g'�p��$�i��MU";;\�r���^<ʝ����>�U�F�y(�ݻQ$���H%��Ϥ�.���UԏY��a�^Qa����/1�0���(�t
�,mß�$��Aʎ�p��+�\���Xѣ��zwO3D����]�oB�p���y��o�d���c�����:��az����m�FO�y;I�suɀ'8�7(t��7�f���Dj�GZ�?�}�w���B�bs�B0[�����=���'�-�*�_�U�9�y^t�5 ��H�+Ab�s���jn�jHY?���h$��Љ����ٷ�=S)�49��V� PU���dwX�p,�J����G`�8ݽ�$%���[~N�^91��q�{Μ&*в�9Ȑ_�jW}&Ypx��/��>��]!��v�p��07L�Nmc��`�/�/(��nbp8��.��2�dN��PQ�A������G�۞��]�QUx���FV�>'QpDb��Ȟ@�������8����QJ_���GCa�8��C�����Ż��7a���w�o�(��Ȣ��?�P ���(�fm)U;�̀��X�˹tL$L3;N�'R���?�R7YO�Z
tǪ�*Qz�u$*�5�gC�k`���r�e؝������-�P�I���DE���G� � 	)ȌP<ۻ�N���^�`#�U�J_��K/]߉(�~���?(D8��AQ �`���E%��|��lT׺'����ۍ3t��`�8�����.f���a1�l@h��S���$��-�a��>������t�B��~I�ȓ/]s��S��*ɟ���t��t���>��w�F��ޙ�ohP�g��S9��1P.��u��[�P�Qv�5���cf$X��4����T�Lfd�l�u������ƭp���KӅF�x a��g�#ҷ"S�F&i-�o4fD�X�4�����g�'��^�}`<�k�K�g[�����w�ɸQ_�]�<nfg>�4LҀ�Uh!}��X֡��ߘ�~q�F��r5�vR�3�3^�]q�2\��TR���0whG�ۘ�1���9Qe}\�x�}q��{��H}'/��	Mf��WÖ?t����1�� |�~�@)�OV-|V��}�E�^K�uY����孀������)Ћ�[xML~tC��s�li  ��@�7p���ꕷ5Y�Iȟ~�|^� !͂��8 ���`��$��J��ͻx��6��P�=#wTp�>L#U�����c�Mj�,F�o>\��ē�j��v ��� ��^?��9c���I3�x�`�Y���bLX���Š�V�Q��3�#<js�S�`1���g�wa�![~���Nװoc������:ܐϰ.oozT�|�fs�W�{8>4��Hr�Q:<�/���j=ZI��4�L8��-��@d�E�e���I��Mm�M�5,�M%1�)��7C��������K+�]����RX�����A�D���[�=��$Y�s������%O+_uĽz~{7���8]�n���r�Q�c�0F\a�C�4;?����˺W���=�C�d��O�0���e���<�� �d�]��+�)G���4��˟��b��u�3���q7�� �
�X�&SֶH�՗n�l�� hK9�슒��)�t����H�i�����W�� �a��t�f�yQn�m��nEr��T��i��S���n;)���q�w���|��ݑu}�
��!V����
 �N�x��#�S&��n�nR�-G�N���F��jre���EǠ�z�Pl���K�z�:Q}6gj0K`]~�8*�[�{��,}��X��)��u-zؽF�c6},�1�Ϧ����}�`9 ����� `2��cC��u�m���o,�#tzCm����UN�i��$Ր�_��� ���B��V�)��,A7�<f��ui� ?��E�+��Cl9��ܩ���8�66����4xĎ���Y^Z]U����?��X΍���I��ǈ��Ϭh[��+	����]r���\��D4����?S�u	����|\? ~� �T$ܾƛ)�����R(ԀJO��C29���&LB�$D8�?EN�p���>�턕[L�a�w��7|xAJ&�F�b'j/�,z*�L�l���g"� 
ÂϮ�eȔ=Md8�V��Dk�As�R���w�����`sJ�DԨTO�G���p�q7\�3�-�\~����F�=)Vָ�� ��	�<W��7ڮ+���Mr�ݛ����ź�1h�^�M�t�2M��F4m�Z�Pa����D���S�Bնww]�lq���ۃ�ǉ���O�ҕ�6{5�w�F���f^��mUYw�D	i���H�w|���1������Px3e����6��W���²���uE�����¦�M�R��($hM9���!O��A��@ZQ�b���͡\��*٥�]y�I����sC�D;N(���@R�0�(л�փ"(�TÅ�%-q?�만ZEo��
�-��A[�kh�ף�;%�FU��Y��/J7��̈�TU�ʋ�����u�d]�?��p�/ H�?�@�p�2����RO@l�@�aV!�ݓdv�!`�کָ���H�B0�� �7T�k���_�ܰ���$�Yx|*��7�:�����{����t��M���������Hט1�Nz-I`8H`w���h�N�mrx��e�rW�����+�{�:�DR��seQ���0��8�%=�&!k��p"�W��ة�]�� g�~ُ��`��(߽��k�%�j�2�6ɴ5x$��}�ߩ��X�X���-$�e�|o�?5 ���3B#�����m�*.q�u@��GF�jH�H�N�����}$"��>Pִ%�m��?�֭���z�˞�G��V"EO�pu��� �{k�VU*8���Ү��.�GY�"��#.Vi����S^&���1O'����]���ٟe>�AI��6��ZI�_>Cl/|_���[^,�~Y@� ��aO=N�Pev�j�v���,y�_{����õVz�k R;�ֽ��Z^�2��_ �x꠺#�q�A>���Y�j�`sC5P�WSUvp�89��&��cR������kxE]U�A�.��Ń��e�P
_h����;�6��a �!��(t 9V��>ȥ�"����b�C�
5_�.^U��Ւ�n�
����3���	u�.M;0�{���āG�UR�b��|s��+*�O�eE��!�v>Sp�� ��BG��o3���v�՛�1��q��6l�5?��%�"��a��+�br6�65H�p��#`˚	����_�^�Y�kV�,	]u�w֞�c��~�2� ;*m��Y�5�����Z�s�wTR�%qZq<C�aD'݄i����ȅF$O�Z����97|����+˳����\.�1 P���H�^�q,���=���lL	*�WmF:p��~2�����JS���#�� ޴��ݸ�X0��Y��,.�	��^K�f��4[\�9\�	ɷ��5��LLU.h�͍ڪ���e�*9d�C$Ŕ��D�S��9p�iSH���%Z�Q������z��*�vdW狕���B!YI-h���M9�d��e��r|���λ�Ys.��n���"�/�xÇ�l�;����op�
�-~�j��ol��K%v�, �֐�� ����nD��u�$+4�(����;�N]�ޥ�,��X��h!�F��� ��9 w2�	ؑ�����fs�K� �Q����>s�Y5P�CmG\E�
4C����ّBK��w�į"ǖ�ή��n����C4��8̐��e��S���<���uJ	�3���ߒ��6Y�&��^�86YsH(Y�{� E6��d�@���|u8��lbw�˃���W!�FM=�������Wx2�����^zO�G�&(�������u��g���X޷a�?���N������'��<<,i��-tR��e���b�?�9uz O��e�  	����m�;��.��^SxG'7z~_�]��wb�|��-_�@�{�RN�eL:�t�wh����p��OU�*�o�]n��օu;� n'+.�|j%���<���:=Nـ��[Cu�cM��b��WJn�SD�3�*�}~�O�Yĵ�f-����f1#MY�J"rotᵂC;+?7����V�1~-��*<$E���S���aS��5I�
���]5$��VHNDUq�
�?���$Zs�'ɯ'>���C�y�N���J��+>#!�/�q��F��T[,�µ;B[h�%:j���-���%�ť�Р����o�V�(uU��HNK<
���rd���䮾��gL�_�L�^�K��ŷ��q�I�5q��l�F�!Y���s0s��Ҥ�.��OQd���.O�?�8�hf�v�s�-�����
���͘ Kj�x�#JQ�QbC����h�Vď�ڨ80�2*:��ʅs=@aM/\!j+�~0;���+�FzW�҃b������0X�wz��q�"5��LLД����0��^����������{��/�����DJ�%�򆯞C�rx�RR����^@���T������x|�5.�=�!�c:���s\�j���5U��йvX��3R�g���>��f��^^ �`��Ц���U��7�G�*S6�86[:��2<,�8o�#h���9���y�L��O}kt�H;x�~k�'*X<��_�������&�M+�n	��?~��d'�B��^��ynB�ԝX,���kT�	N+��[wժ���D3z�)�x�	��-3���w�C:�,��0�Vu�uܑ�Lg�����s�x�HwQ��V7��
�����'�x��ɤ�ˋ��J����K��鯦uV�v��F���G ���'���G�9��U�]KL�d�`���$0�:���� ��ˀ��aN��OL(��T��3���8Bf"��4�`5&}S�����v��o��R+��$X�}1��Pr�*��jh�*o���1z��C%�*ys]Dp�u&8d��!�Ѩ2�����FF2x&�`���C���o����qd�dv����V7�%�x.4��oY�D��
�w���iP�`Ջ~������Z����A�5���I��˒أ�)SU�T�_(�0�I4�J��Dh���h|����S��D�{�5�0�0q�ٹ�6�m&f�[�B�ٔz�S�]jZL�ߩ6�̱j?ԧW'y3ʇ��i홠����H���do� ju!m��"no]d7r&�
H�<�,q^�qN�EL`�g���L�6�m�8/���,:�O��+���9*��}g�=Rn$?_�{Q�R2�Og��M�Y�'o>�w�6 h����sY�D}[ʻ�2���0���k��ٞ�a`��h��EJn<�KV�<��<��I�HZ��U��b��UGC�Um��rL�r	�\����HI��Bq�rwG 3'�R9[�׀�(mt5h#1]�n�J�A^����'iC������,O~�����և��J�t��}n)���&� j
�_�SV��ʞqg���|?Y�;of_��������%�!�v�D=֛�{���C_�i���������UY���L$��b���.��u��@��82e|%%0��5h�>#Ejg ݺt��/����������M�줅�2��
[����L�O<������ڟQ�-��^ 
mW�&�w2�#(�m����x8�X�#�G� �h��X�5�^�UaQ�/�C��s��0��~*���om���</�9 ��1�7�E&����*Qt�'��Xag�5��'�rLW\�/���mD� ��i#�o��8�/H{�Y>I�`4ơ�'��*�`����Z~OY�A�vn�����6s>H� 	��!W/R2`OPk�F������e��M��y�g�ǹ�{�����lZQ��#�el�a(����o
��6^G�����m�q�e���!���>�m'�}�W���{
�a�:d2ʪ"dc�4|5�&�!�K�{��͛��V�N����MO���Jm�cu҂���^�&&�L��P�:8ﳑY|p�����W�{,'��C@�9o�&��}x�����}R�������G��VF�����v�j��R�G�Lu�4���gJ�v[\�v�ȁ�/t2�8ү�џ�]�2�nI���כZ��yN�h��s�߬���	� �o^t,>*R/��[�@p�x;(�0j_�V�DJgZ�ͮ}m#,���5bO�Ԟ0�?S���L,�.�C/����b0 �g�+�*�og�N�i�D[̳p���4 �����&K��������jJ��6�0ع����+2�D��h��L�M����jWA'��F����T9��E]��O�/_��iP>���Zg~��i Ī����2�nY������#�[;{~�s�B���~U �9q[e��4��xc�B�����������=q^�Ddӌ�����J}
?��_ ����n�X����y����d6�;>�s-�H9��&3q�e�F�o��a��@��aﺚ���C������(�VBqn�d�>�8�#�c�R�7�RP�Ȕ��`ŭ����ҁrJ������;�����k3���,����M��$���jU�����w�{��s`���̊Hzy~n����	��9=�%z���ٚ�{��]M��vfx�]b�>.rg
�FecZ҅/���E{�n��Z��ZWͶ!-���;*��l�)��F�=�h��Z6��$�e����t
AA8����]�1�� kwP�^�{�͚0#^j&�� rI�D��#{�C#����GW�<e.��V=���1N���j����� a�d��5�����f�gH��rJ��q�ؖ͟κF+&�R�dE��ST�2(��U.H�"螉�սJ�r38!�ʢ����4�{� �*��qV%@e*=��`-�DQ�bA����1%�UT��P�euo��ɓ��n[����ݣ_<��D�� $�\�kYi���>�"��3�Y���^C{��2��!
��8@}v�V��4�L,;$��dߋ�`U��*o~dn��>f�?3�RKʛ�Xg
�+M,�XY�)֮�`��'���^�w��m0ȅ5�=4-|L�Q��5|)T�9{ձ9���{���hܯ	��*�c�D��dv�����M��.�Wiw4��,eU��~���Z����=�ҳ��< �����i����ª�8����܁�	w+�&�li������x@]`�Aɮ�8U�ϡ�<�f��"�g<'b�" >����j=#'�{��ǟ��?R�2p�I���r��E$7��3��8R��[�{�A)��x� ��8.+���-�`o��v}حMG��]���p���E!�*�w�Z�9ݮ��Ov��.��� DN���N�W�.��O9��F�0��2$k���PtR$�$�[ص0�ji��FYS^a4%�	�����T3[|�`��vV��b�`W���ڳ!��{r��T��.�U�l��&ݻ�ƛ�P��ޗ���p�P��C~��#Tt��9�$V��8R�o�S^��[�{{_&�S����VQ�U�P}����Yc�N��j0�-S �}�*������?�x#��	).ZRC����E�A�#_;�Vg��'��=�d�/{����aR9�W�B���fpX}9"��"vF.�'�sc�Һ[�E�vދ�hvz�jv�p�cX����cL
m�(Po&P�֐�2fw���+��h
|:�fy���YdV��n���B3����1�t�	l-B|B���u��"��hVM�~:����Liu�ϧ�R��<���}����(8U�/�[�l]$��W�R�r�~�D������(Æ�i���8�]���S�5�"F�M���s9N�_|�I�c9�ZS9l�!���59��@W���ę��[-�/v��%_�.��}�܏Dw�,����.gC7{��_��"�J3bf�z��6��]�����SB���'�G�OM;;�9�=�b��F�4��*�	�g[�*�9x�h���R��<(UMtm|�8%�C�,ViC�5�t&i���Ѥ���A)�a97�
��3Tᶕ�d�T�ޚ%oO���Nݙ�]�_��*A�@ 
!��t�_3	�
�I����u���}'I�����"A
d�l��e6�ֶ_~�i��٤���$�\��9����
�As���YG~���mƲW�9:v�/�x�@����Fz���;�Z����|�{����g��ǖ����C���d��6d��r.�*�!�Q=PuC��oC�4t �>sf�J�=D�WK%y���{��)�}"q��1mOZ�w;)�.�Ҍ]��x��4�Zl�k�����v¡��5L���"�|��9�4U�U¥��$�{���U�kuZy��=�f��:Y�����~!H�N
����Zv�TbT� 9\�h�^���]����p��L����u�;��Ok0}�=Z�ї~"iB_�����>M�&
����lF���w������+�aa�k��B��mw@�,�ʧ{�v���~g��9���Z�!��[���p+�|CT�ɔ���+Od�53�������򔔍8O���5nm=y�s(�'�{@���[:P����ᓣ'ɍ���#iT�	� �tܑ$��ႃ��sR���ǣ�*� ��!����C��H��c�jy�_>�hAJ��~Q}'��2��r����7���į�޾=IB�;R2��?��%�Ƈ�5������s�>{�������V9u�#C	/9�Wb@w� �	����Jr�L["�O���2�ȝ�O�v����rk�`���X3�2�2�+������k��p��J�2�&�(���a����!��{����jb��~D���U=L�qO�7���zA�
5�\����F�2�̤�\�0n�?,��Y�t��+ǘE�� �ն��.�zF/�y��[�?��Da��{ǉ�o���p���R��]➫��ȏI���qe��<�,���
-S�ͮ���d�}��WQ�����)�I=O�-�h���ä�kK��_i��ͼq}g+�v��7,�+=>���O卓M�������dߍ��>>88��4�sMf\���˕�<eS*�����t�olL]�3ݬ��鸕�z���k�=(�ې�_�~چ;N�K��g���$8L��O.:�?��6!��	���o���5 �����{_�TR�o�M�ݸ�-�ǃ�v��-^�3�n��E@[ǘP7�a[@��)֩}Am|�і�B�f�[��B��g�}��:ݘͰU	�jd!�6`%�0?��	��~�")���5��TW�U8 �ݵ�l��N������*<cH��*��p`�9�� _��0ϗ�	@���%��U|.a�P+�"ӣ�ɒXj�n�ǎ«������RY^����س~�p���.s��"|�����5�&��C)-��_��K��Y�l��I�2�Stg��{COӿ�Xp�!�i��)u�[KU_�E^:��XA�
`�0^ n�|$J��r��G�B�B�����R�t@�M]�Γ���w0?�n�k�.H���9ZVl}�!��~s1�ì�La��b�-��Yω��6�x[oGy�'}6�߮Q+k�X�#8��#B���>F�VN]��/��.z�P��eX8�Ϧo+���"V%�ƨ54j+�h��nޤ����q3���Q_�U�d_�e���)�x B�[�Ë]�~��.�����nS�!:��F:���@$ԟ �6I.G�/A��&�x�8����[���Mv�hJ���ӷ�m���7w�v@q���lT�6Yt���@mx!UN��o~6*(�V&]��� \�Cɐ>_p-��\��U�Q�9�w*,��O��z�>�\���t��,2����u�g�����maz V]��Ey�4TV��?�ݸX9���L�v�gYweO�������$�zoM&�d������Fq��b1<T$��~g2����(���i�>�6��
�kΗ���2��=��T4�P����m`z��>{�LV%<1�m���m�BW�[�"Z��G�d�V�>��If&:BuS��*@�+�09� �M�1����!���}�m��/�~���2Բ$�-e��ցD02l�E�Jm�@�}�������s:��~��]�x�G�sH��AA0�6rAey�2��M��⤗��f���J����8m�w��0E�#�HV�?b��=`�_d��;>�#[��p+�ۥ�ܜ�^�M,bٮ��H;[�P�1�7�#��������5�@���ψ�ܠuq�H:��
kGu�u�عya5�6���z�{ s{D�DH@WC(���w?����p�^�]��=v�܁���흡u�%�NMfi	�t�}
v��n��3V�Nߥ�ޚ�,�kԥ�#P�ߝ�2M��	��0�n}_���ʹ�nR��D���(�-~��(�r����>=�? �<Iw�c�^-_����+4ЮS]��7$!U&�{R�D�>�0Ap	�#�����7� �k��PĬ��T�L�,	��b�t�AG��ä{�ai͢?WOQԳ�F�du������wL��ۂc�O+�)@s>��ygi����� *l�XJ3�ǡ�f *�P��f�k[�7G��w*'���x{�<�-���Ψ!�c
С��h�Ч[�q�O@�ރ!0�/��z�e�����7Y�U�(K8�&�g�^�$}��SŔ����2G��!( bwɷ�!p�{����)񐠴��m/I#	�l�5��M�f��~�L�|��%շ��w?��w��&\4�-4�b�#� �2��.�Ȱ�W��D��skF6��p���!��r�c���[�>��I�G��T�>���d�l(	c)��2Ik�.�G�6m�Nܶ�P��lSpj��@�n̳1#j��GM]�O�����u{w�Y�45�d�rJ>�5����J�����/���w쵩�t�b�=��@
]�V{f�Y�%�'���3`�>�}��L������ ��0��i�C�k	5C�Յ6y)9�U@��'x�"@�dq�[���\��5Y��5:Z V�W5nb��{��S�����Qe�����,/f^���R�Q*C̴L��p� �Z�P�Gֻ�qP6.�E�W�}��������2E�j
c{\��i�$�M��n�i�|g�O�����A�7�-^�TDz�7LPd��JY*N����R��L;O�̓B[�.4!�������Yp�43�r�p3,�Zm'��A��1jsh�ۡ��'Ѐ�0�y}~�s���dK(���֬/ҩ6�Hp=��?$l�|y�-,��U�w��~Z��Y����&mGC��i�<�o�;�e�J�H���=K����R��āO�PuMg��?.~h;�aO�v\6i�8�|�K�����3��h�Ni��,�(�S�)|����1����� s_�h�c4﬽�+ګ_\17�����T����9�R[��:�c�࣯5��KmV���� ��^�hb�Wg�JSpP �Kn:�̸�,�"��� �1�5���h+QTz7o9)�	�%(�QĀ'~��X����k���j+����&��=A��x0�W�����Ǚ���3O�Z�K��(�d�Z��,��w��n�=��-Y5^�h�L��'�m�V|G~�B��v�����7����K��v0�p��m�3�������Ϝ8%��U s��'��&�C'⏚��Wp�K4�0��*L70v�lt��WCl#��	Sr���3�v^�g��HT"�zP��9�'�f���Pʡ��V��_����ċ,�7���CmW�
czg���l����TN�kj�l�} ����(L�<���&�_����H�u���Tj�}��/��������7OB9U��{�Q�^ɺH=�A��h�x�9S�M��慯�[�ة %���)����zh������ѭ��o�@p��Y�s��������h�1�Y��-#�,(��p*!�"�$:E����[ d��=�?i)��� աE6�P�@��M��j;���/�KW���>Oś��_�x+������\l��J�4�~�߁1����`7�^F��9)t����GrX����Pl����
Bɗ\�M�C��^c�R%z{���0a�Bt���(�`�
��pՉW���1��;���ڧ�-���[�g'iw��X^��%Ħ��15��v�:�{�������@K�럵����n���J��a�9y���4�N�C� �S`�<�t�U�b�E��$�e��(�j��Jq̈́c:jG�T�^�{G�K0��h�or�͖�����m��!戀��ugnjذxĿ?������V��_<x!n��������"�N#��t����EpR>�x.�	��j��+�m/k��f��g�������Ĥ�׾e�IW�%p,L����>LQ�v�d��l��m����R��!�a�r����X`3��x�0����:�����ꅈ��fIA��L#�X�B��+l�Oo�~��|�S��+������r%;ŉٚ'��N�F~)t�fc
�(�y�!"k]C�I�n_����孡�B�L�U��)aÛ�Z����!Zf�2<�+=��S[�{��������BI�H�Z�\��d��39h��c����(Z��5�j�|��.Q����vp $�!u�r�9	�Z��ުO�0��bT9=qľ�@����$O �d]Z���[#&���EI��4�������R�0ޟ� ϧ�fI��0S{�E��#��rS ��"3&:y,��B��=%ΐ�x3��\�����d�]�O.�JbyZ��A6I�&)hӯ�"*kƨY�@ ���\p!c7�$G��j�Q㇟B��όug��"1��	~	�ʻ�m�}:<]�M=/�.��˖l�������?�o��#��ٝa�e-�0�e/�~~�VN���Aģ�p�d���\�n�uq%��B��`�D��p���.�a�B�Bq��N��m�N�2U,>�4Ŝ��|��g��?���\�;̝E�)c���N�\��[��שjR�]�1�	�rC�ھ�gİ\���dͨ�wBwM�y[
͕�r+=�ޥ�kq�K�gPeޏ�@�� (�(�%߆�uc���>D�2߶Fl8�j5/��9
A��v�oaqe��k��˄޺J�N������◹���N<�ƚ�ZĄ��װO��7�I��
�?c}_*�l)�$B��_�����JE��߽�
U��MB���e�"V�������K?oS;?1�1w�W,��>6�X��x�s2(Jҍ����"�K��g�i���ʣΘ����U	@���P7q��7kc$�+h�ۘ]eŪ�.�����o���T8i�S����UYح��*U/
5a4Y͟���Z+ïi���^5���ڽɇ�˫6�ǹ�F�C
��yzK�Cx®��&<����f�E�fǎ���rr{���s<�V�eu�ĬH"`�w���&l���	�h+?�����͏���lX��V}!-�5���hn�p�e#4	$`cy�n�`F<�_�E�U��'U������*|����w����e=}I�`k@�^��WE!���Lg[Vlt�5�LF�r�E���$��C�JS5���wK���W�<u���JE ��	����W��S"*Y��d��?�u��-����󨂫`�1�*��:PL
I8(W}��F�gLݽ�W����*�1S��g���D�/ό�όԳ���2��T*�^^Ds�H�B�qcQ&:�}��sg�ۚ�,"_�G��7C�R��ª�o������և `�øb��zmqqN�m ��qDFs��}qBX1�\j�>kR	,�����	�]�f�����\��	bE�n��]�+��Z�ꋇ�� Hj֑�se]���ƍ�R�b�d�4�YY[<<|9��_��E�&�q���f��ǒB K�&��w9�O��쥮����]a�Zg�;w��8�2�a+���4�6�z�BP%��A7Q3��0�z��ND���)F����&��?
SYR�<�fΉ�&���3�%��g�N0���e2��$E1�J��۫�d�x�37iRP�������a���H0,L��a�^ $��E�*�\�*wO���5p�G�T}*�gZ��^(5�&�^�[�?��71��?��?�v?f�Q�[5�u;���L��.����v
�{ ���JD�lhW���=a���XZ��OĽ5�΁�����(���� a`��o|�>sۑ$�2�;9���|me�i׋�S��E�4���r�:�+�����PK�3�ʛ!|7� +����e�e@�;�����Z�I�Ԕ����gE!��i�0��V//^�m��/MD��"�����y	�"����6���<����ΪOD�	|өژnK��>�?���--P֩�vk��Vȷ�s�V�0��Κ��=w9P�m��Hj��M�/�����F��rF%xm�.6ړ�Ma�x��Ҵ�r�w{;;��Y���5�"���al[��j�	����b[KݨÇ�}�yq�G�dc�J��<�j�*��vҚv��oQ��"q��cdYJ
ƾ(�"i�gw_OCy�4�'�.x�J;f��d#n���q4��ۮU�d<աP�^��!�Tޒ��T�>lJz#t��Y�o��#��o=�ɮi��&v��f�f�p�6�5ivP�%>Ŝ��(�I�ӿʔ@���Ӝ��9}��z�K_y(�+R5Ԗ���IWcbSu��k�:!��H���7�$�;�%������a�e���Ǔ��) 吟��l��+�{�S���n?+��n��K�BS�]4y��o����$��l�xd�}g��RݍEڿ���r0^X���M8҆��oP��R�s�d2�O�jg׍j���� � 2��ز(�N��Qf$ovbf�1�0!�*h�[����"��B���4J�Ϙ]�0�{M/��QWKP�PΗ�}�����#�79�ѣl��p]�O*��ciL����B�t�q�k��o���-�
|�=��/>�c���_�ю��!PFk�l>�W�.XߜS����×�{��޳���Ӝ>mP7y��mW�ٓ>�'X��o� � ���q%�wu\�Lj�8-�����h"a�ڢt	��0��I�B̲P�-�)��E@H�� ��:���t\\��x=�}���nF�:��������mn;��a�	�VzA�ۇ �M�1�l�w�mWJ"����r~��a�j��q�g�_PTh&�	U��;�2�w0�ٵ�WR6�*�;B�8Xb�W22�h<�¹�S�e5�D�Ys6�R��8�f�OXavݓZ���}q/���|��b��s6?������%x���
n��\
e�{�D�E��/^xZT5ہg���"1���d��d-��&�'�6ա ���84���;\�"��d���P�]�A���?���"d'�SY�r�,��B#�ЪxF'7D,;�z���E27����;z߱�>�ts�@Eө��&_ �B|�!t �q輬G ����K����3�3D0ƙh�k�V�~<���O�
��îT��e�;�k�����4��ӧVg���[ ����)~"��ZL�)I�.@�)qA�����%���t#�2[�����{����"�>,��J�U
�0�RbH�k�Ku7�us�uؘ(n�BTH����(�G����wI�C��l����͈�7.�D��Qh�-}<���W$�8[���D-�R�I#Fs6��XE��4`�<��2A����JAN(H㏫��0$�׀����k��k���7`˰�u�Z�.�g�i�z�!��sr�2+$�C�Zn�G��kn���9�-��
)a��عͰ�H�f�$�+�o�n�W����S�S6T!�*�P����@�C��rHqob���Zr�o��/E)Y��CVt���4fH-�MW�|K$��2M�4�.�iU�ӎQ@;�t��s��ޑ%8,�#~��UeXȅ8�̗4\�oTjG�O!c3�0��8m�xzSit�$[��1ߊf�E�.+VA(���t`� N���r���6���9Y��f�8�j;��PVY�i����M,/�����}E���Z�g�㤑���<���B)%�4|R$���Fcf͸�'�4SP�!m8}�T�o�w�H����i�qF�A�Z���i{��g�)-�w4�KJ��������<<�J�d	*Ma
<T�^�M;Ԡ�lwvpi<.2(��*�֖T�����%ݮ��kZj ��@9�N���,�0^nΖ���6+l�v�Vl���*`��OY@��m���nî�x����t�NR{h��'>�|͂�Q9yw�#���*�H��K�[N �j�`jʒ�����H�Ԙ���K��l����/%hj�H,������S���0�{��A�..�g���{XAH��:�d��sK�]�Ш��1��Ͻo[��������29e���¾{O+U�S�Y'Li����Ĵz�����%�5i���X�h�CW~27�N��V�׋ �[�̐�Z���+�b_Apkz_.J��̒G���'Aδ[��ѵ:ր�9��j���"Gw����Or��.ϦDK�m�+��
"��$��{���[l�)N#�7/k��tu�bP���[�����T莤�e�'�A�1��-;��N#�̐.0������N8A��X�`oM�lH��{����bA�B?�߇.�=%H{یJo���Q�4�l+8�ߑ�Ex"SP����0z�6"s��&��(Y�F�����ew�cc��x�Te��Ot���P�Ө�������OYj���``.LgJ��]M a