��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��0�׾����I�G?4�xC���-����ip����)ױ	J����]d	��$��
��Y��=��A�~��?#���@��:�-�=-��l�Jl�T����?�s:�Z	���-�F�wm��Z�<�����m+	����Y�� �z�+�A� "�R4=��GU [�]�:#�Vφ4�Ik�������>xG�>E���a$�Z�=hw�����¥��_n���Qی�
u,*L-�UQ��ʛ�#�A�gըO���R���~�!,t=���j�3l����
5N�7�!��q7���O�s0u7X&3k�T|�2�/�W��;��*�c����@�Vg�w� �Dʤΰx��!x����:p��@��[t;�@�.���M�%R"�Bu�6���zSc��*���1���wk��c�SJ���I6�f�!���ā�0��0vIz1��yg)>
v-�]�.a������`�`�5���1�Qw��|��'Z���^�Ԥ�1�W�R�"F�3R^�y7��|�tp���k��d���=|3:�n��Wb�����>C`^����鎶�L��n�T����W����94�06���G�'Gy�#FF�B�z��a�2�(��"~��E�{x�L��=,�Ƀ�S"��&c�c��ɤ���N�Y�	?.��lڈP�� GST�]�?����õB���`-�i�M9�uK��V��F��v������]��p����5��O��M���>�H�.��5$����:-���͓���w�EU#�Q���$�k����V/lE]�N 
�F�<�[�؆�P(���!M��\ǒo�+����(��*
�3'[�^7K��#�Z����P�{<rޭr�Į$bP�)�ʼ
2�9�I#������y���Y�˽`J����2�7�����D��KPL@~��k��QDM��g�q�m�'�L"q����/QM}&�R�"@%O
+N6ӤλOҔ�n�������vU��tɗmz�̅�]I�-ƽ��֗mo<攕9>(�}x�jG�kc+��	[�[M,L��MC��L��5��b9xpUy��ԥ����=F�+�z��wZ����bU#��b�8d&�?�"0��[z�]J#�>�V�0�z�l���/
j�c�A8s���<�1ӒPJ��|W��+c����O��!�Dp
G��M��O�:� 2/��B��&.�N�}},ܝu,���,W0�|%É'�ѵ$��A���6�כ�w��m�&I���
]gK�RJ���u�X1�U�ﮇ>L�e��-(�L��w�g�Bܧ-KT�vV��,��Sd��ݵr3��Lx"�ć��M�x�/��_�F dJ�pk�f�S&@�*֮�vk�5���)0�����4?�2�{��� �C���e�	�F�ʆ�I(�ā���dn�;�#:f	|u��q��$��*��"��&��I�;$�cȬ��$�af�6Lk�w���`B,SBPM���~S��$m�N��~�����!*���C�6e���,��x�!=6���k���g7n���2��Eޟݨ�&	o��]{�5�J��yAㆄ;E A��� �I]����t�9���Uh��vme�� .���O-\���}ЧG&�髅�{G�jE����h����Z���پKˬĶ��90�SK[��x1���z�hأ�,����A/�Q��X��f�i}�<,Ƕh�_�X�$M��g�Į���E�/�ߘ�Cn�4�_��Pn� 0�F�Mt.b�F�3�:��db
V��l�w
d�M��M4[�;%m���0�J����=5�`G#�����(�k��dIPc�a��ݒ$�u�*/�&mu�}8�jQH�FF/�7���� uj�+f_�I��<�e���2//��U�`@Z4�ŗ�Z�ݦ�����4׫,�:��{�6�j�lg�����
���Rh��R
=�5�_�4�3�G�n�*��gа�XHA��B�Y8=���4z	4�ïo�v����_Ue���c3�c �`\:g'X��J��_�m���r�����u�!.+ W{��eHL�~P�'�0�ȳzX2�t��A5��(�b��&.����>D2���gy�`�(�w�����n��M�����-�S�8P~�� 4��<���t�$��żs���P,5'�)��"�[31q���� �D����6ha�S6�p>������3���7Dڄ	�	u�%'1=YB���N����,�G:��/w��[F-��̅;�w)�n��� \��]�Z�����MeOR�(���ޫ��oU��ڨb���#�u9�8F�C�6Ř���đ�`o����Y�v� .�vAx�>�H�t"Xh��>��G�e,�e�,���Ō��y�?��:�C@�s)y<�#G����S�ޫ[S`�B�� _}�O�q���⤌�����O>��Toh�ג�O�Ѿ�Awe���/B�]���<�AT��� VR�ͪ$��`<�%���ޫ���pyP/��̈́_�ϴ(B!\}���"ZM13|O����HM�'-��~x�X�5`R���K�x�����*��zJv[Uj���(V�K����s�J��<��<:yR==�D�ܑ����t䦉�����#�d�kD3��]�g�K������ld�Z����4�H:��,!t�[�H`�m� ��#1�ԙ�U�ڎkW�s��r�I����}s������=@��+��9~Ȥ?��g�2�*V�1=(��=�Ф9�=�y�O	���>�����S;�Dҭ5H���:5\*�����+�	�k*ғ �BG���q��@p�bsR�@4�`�������W�0y���<J�q0j��cfP$Ϝ�X��6���+����a�0�zߒ����yy(uLBJ_9��5���ԙ�EJɲ��U"�XѧP���1m
wE��goˇ�d.\ �����?e1z�H@��v�TC�� K�ڿ��U��C݅6���^uN�y�i�ph���߅�}pb�x���D��GP���iM���:��rM���6��ZI��ýVQ�2���=A��B�t7,W�F��|�qH��:2K���H+�\�+@����Z��}p�iQN���B3���m����S��u:S�]�2?9y�L�����;��شF�������{i���x�Y/�_O���`�2�*�Y�t����Q���Q��=\��&���J�����/�'.�L����ﷀ�EO��l���ڳcY�/1& (/�bl�X�� CNhH}�����.,�P9?'Yԡ:Ê�P�Z�B3��$=��
���,:�v���4}	�Nb|�[���"�����N��� 5g��*I��a��������4,����'�O�]��3��XL�	Cմ� 2U��w�q_����O�:�ڄe�N�,m��@)���t���+e\���*���� ��@�jID�wʯƪM����eƶފڟ�Z�;��f��/��S��k-�P�9G��ï���(G�%�	X�p�8��H�*A�]$[�0�a~��ԗ.��ͪ�W�!xq������m�2�нݗOK�2����'Ag�]�
�&��1w"�LR�>{s�k�����'�ɬ��I�mM^x���M0�4	$��q��Mlme½2KZ�	G\oؾG�������>L�͸����(�)�ϕ)��qiYE�ތ2}�H?��:��� e�+�JX���&7['aɌ�6��ޟ��g��QvZ�� ��W��OI1���z��P�HR"Xo3�D{jJ o"h'���N����:)��i�����P)q"�DgC�֐|
�C^k����ڳ�8f��S���R<���O� ����%�x�y�46�Lȷ�ޅ=�#�E��4n�y����4��2�Oe���?,L���E}B��d
g�)���t}k�4Y\�W�1d��	��}^�zB��_����<j����<�p��,UqnC_݉�����5����L~R�͆�3dR�%ᖁ��i��Q���'E�¶}��9:�=�����Ԓ��@�9���(�!��'`�����D�,t)�(X�
 �'�0�4*�Zg����X����w�~�#��Ѣ�����(�gz���e�M	ʧ�O�9�$M��h;CG�"�u�d�����h���f'8�&�\�.%'}Ŝ�g-!uL~ RX�h��G�Iص��n�����)������&Ѿ~	����8%O�kJ.2��#䪶 �Ů�R����+j�,rO��a�����w�v�J��ⷮ̐P�J��Π�Н�>�"ޚ9��H����UN{��HX=s����l9Kxɼ�2���C�"������+}�g8�����lQ�A��ʽS�MCE��T���
;��U�0Ȧt�B���p\�32�Y"4���wS�Ŕ��͜Q<
��t�Ӡ��!����&o�~����&"�3N����Ѫ���Zs�Q(w�Y<� ���,�l��&�kF��]�^��L]B�&k�]GcMM�}�]&�c͵f@FH�3O���}�!R�t��\�s+�I��!��PD�q��i������v�4)Ҍ�ܖ3x�I�ZL�De-<( �J�����/���ўAF_�.ڏ���}2`W�q"�YM�[�4�(�@	M;k��k�5q��>
%	�������i��Ä0 T��K��a�&ڋ�׾Z�Z��f�6g��Cs�Js���US��h�V� ���� d�i]YI$W���qҔt>�h������Qr3,n�q�j��q���k�p[L�&N��7�&�� S�N�����e&fLe~b���l����̀�� Ҁs��b�^jKP(��][���������ƈ�)������[��8��/q�)`>n���= \��H�5ߗ����H%8o��sV�ZƱ�0&No���[Dkhv5���f`�j�ɰo�I#/[Ut����
�4�Jn��ܤ��5��qB�|x$Z_�_�2qX8�s����OK�d�E�ҥ��8�Z�t��K�!<��|�g�<R#.��B��`�ٽC�6-ڴ��T4Q�?����Δ&�*�ꐗ���(��4����w�>K�M�CBB��K��h��o�?�7���8W�mR�s���Y��*�E+���/��9i����Rq&?%񷞧Rۊ�?>NoTN�Ƒ4"�	�Q�X����0�$a��=�Y�y�G�'�8G0s͘��$�Kl�i�^��T�g��_��d���9��XZıMPd r��~�Q�|*Y���3Q���/���j�@�#r��Tٵ�Q��C����<�����rj��c-,X*}��� 1Q]������`�u�uyy_�%��x#��'�U]s�-
b�������Р�Y����Yո��%>��#N�����p���	V�矩���M����Ʀ����󂴇���b�_ڦ���8sڬIW�!�v��4���H�����4$*N]��iu5�2@_���U�:0c��/�_���'&��H�-4Q{%�bG�>!ݎʝ���7(�*�v�/�wW4>DY�ĺ#��_$��k�%l,iڢ+�A�����_�M�?�p�]Aז���<�M���a���e���S���mZ��.F�!�T�� }�~����P���j���z�i\<�%<��(j/]�U����i!M�}�=r�\�$��\]�.4��r$����IԴݖR
�5E��K�Z�%��i[6�! �
p"륔�s�W�5OX��Qsi��3��'F �T]���(3�	������AWA� �qX��R< �7fAs��.�Z��p�
��R��l�³B���Z��}t��[��WR�<��Qmx��sp�!1O ���a�fBP|�
hjHx�|i~�Q�!�P�م�Z�@��?��@���/�T2"�X�1>��Jac�f��a�w?Ç���T���ї6 &u���1�o5;�I\�g��l��P�z�,��s��CH�hD���ǹ*`_���e�(>���'ꘉW`��GO��UN�[d��:��=��ͰFO����[�q�I&��%�N�V�УK�S.���/���D�8F*pRBh��Yq��6�Œ��[t�aW��1��/�ѵ	' ��7��S�
`^'�ԭ����"v�:��.������:�p�{��xQR�i�
�(�.��������J��9y���\[mN�Mc�@��w�G*gQX���"Fh]�������+������z+5prW�� ����θq�W�7��}�}!��^#�/�v�	�% _Z�7R�^L8�����a7�E��H�1"�7KA�Co4l
(S�>��DP�=��j�����n�'� ؗ=�)�7r�Ao��� 07tGQd�t����'#\����:l��P������0ȷ�̙���zD~Ph�˼G��*%���l[�5��*a��i`�Ƴ�~�'�%�zP�ޫ��2אNr9�ʺaΡױZ���G�x�?����L�_}>R�
�'5���.H<���J�u�F��v���J@�Ǹ�$�\C���%%���+e�L��j���z�(t�5��4�x��_"�5�u2ب��Z�ۋ�����A���/�r9
��zʻ�� �:sm"�t�g?���/�w�55ܮڜ�֌�[���b*6�$��S�_������n���Y��Etn�N��PF6�����cS�<�x�����xb~b%
w�E��p�R��h]���Y�C${![Y+C=�������{#RC���eU]�y�^o�L�>c�B��-�Xj^a�tyN;���E�|b�f�_r�\�V�Ȱ;@Ge�z+��CnP.�� �
�gb�!%;��n��
P+"����F`�M�9�L�5���PL�.���nbyqo0Us&8��������~[av��lړ��F�G�_1�0�ֶ�Sn'֦Y<��w��ܙs��
ܦϞs�vD��hH9�Pʰb5��4��S5N���<y ��4�ࣆ�%��膗���+E�c;�`<�~|ʩ��p�+��	>���dt�� �g~9�&nxm�_PK^B��WCz���l��'؝Ou�
s��P9�66�HO_�u��B�!x ա���3)�:`�*����0O�ˢ��ʳ5lJM�f�~��O��+�-\��g��r?@�Q�ܠ~���=�o�e_P[��+3��(M>��~�K�ߑ��pD
�CD�,�y@N���~���@o�
&��
7 ��K)x�֟�ڲ���<�a}�
�9�C�#	 ��y(e�)�;�&��Y��)��>iSAwIZ"���.$l�h�uo(}�Hvlj^�y~����S��S���QT{���F�Ck���	OL��¨��T�,d���𨑡�������[���۞N�-���o��ae�	}؛
�"���R+{ ��J{���$���7V;|��53;墽^�R ��v-���m%O�9/V\�6%1����Z�:��<�ئ5�� ��{Y�V؜LZݻɹ3��cVF#��/sQ�E;Zg��*�J�JA�%�[Hg�+�G�&)�ݗ⫺� �������Z��
\zy�Do�n셌C�������ف��؞l�a�pD��|�gLƆ��0a�<�UE`�Uo��Qp7����̶�����U��"ĸ<R{RUUi/�>٤09��4.`����a��b����ҦX��30����~��TUjZ��,��`#�2$���F�p���９ϸX(�
�ʊ)�|wy9q2��@�,�" ��S�o����h�zn!o��B�]	4�m��I�3��l�:�Bd��*�U\�!���� Nob0��8	�' Wg�ܲ���]�iVV�c[NTL!����_«Vf�vm��5���5kJR�2]�4�ߍ�=��3��~`Bs���a�-�W̚Wq��c���*��K��A��nc��VU#} ����D'���hZ� �h���<��Nz��
�PCB��^�Y˿�y���\qϱ]�c�ׁr��c��s��R#*	�~��z�-�M耳��c��v[+�-��H
K�8q���ՙ"�h9�TnA�\QY�d� �Tt��yq.�J�X�q�/:a����VtV�XF"������	-��z/N�Y�O ����i<�ZrH���@i;9L��v�|f�>)8`����u]�M�׳�d �Bc,y�r}��� }`���?�h�W!js)c��?L8j�@d4�ɔS�Vz�l�=?Z�]��Z"�(2�y���#�Y��Z�j����֘�'8�>�a
��Hy��)�p��
���rg܆wV�Ώ�U$��gY=���_��º����@�V��t�Un���+���q��~��Zo�ɴ ��#qb<f��
�!���dxG�����<�+n���$�кc����SH.����Lsa<�<�!ן��j5Ҏ�z����+�H���3AJy�O���ڟA��=a��G�T>"��%U�~��)�3�Y�Y�6�!�b�+�Y�'HL���}��N�k^dUy�s��LLJ�<!��Tq'E;sj�4��V�ޱoW���x���8�	8����Z��Nctib�8c9G����_��m��7�E��Hq��\d_^3���C�2�._���u��7K]YlUn%��c�����$�pg��99�мV��K�K󽆖Ɲ�?�e����8�xp�`�t�����ו��^-?�$�����2V\����w#}=`�����p��g��&�6o��u�&�i3���&.C�'�H{��nJ�I�xH�cK?]B`G����E�*8x�".ゎ�K�B���
���|��z�;UI��I��j�N��*0��7����vKG�g�~�ݟ�eg�j�n�GW���Jmg��2,䏓ɽ� ��h�l�v(��F�&5~�O"Y�g��l��G�[0!G7��$s��b�D�d�'g����D.��lyђ�/��~���u����2�mDjL؀��#�n8�%���FrQ*W�j�(�䥗�Z�TU���ؓ���T�}�D������e\��\��+�Y1x�|s4wq+������8��j��������l���E�MT(1k�hós3��4t�d�&�P�0ctz\1�b�࿣ET,B-I=���O���loS�:��z@(��+�헇�r�N_/,�����ކ��fK��&3��3T�=�R�zЊ��s��؃�	��J��Ƃ���|��N-L4��&1�������K0���0}q�I���������C��RQ��%��ה��Pm�\�jT�0���0qL"ƑY\�s�?�&�y�Q<�ShB���a��3��^��b������Y�?�t���#|���D�`�� �KJu�����:�Mv�?:�����z���=���E�Fu�E/���N��7��s�4bA��FI��:U��v-�3�s�vЄ��"cԘ����S^]�0*����=D� ��}Z�i�	L�G�s��ď?��ű�Ԥ�)�|���"@�\����J�͵$��

xl���z��ſ�&C%!^"ڿR�S'.(G��ޞj��-��u��p��y�FI��d�N��^xߠ�Y
,6�\����FZ�;d�+�:�`�1w�u��ײ�UZ,F���eB��1�H��!�t�K���Y���c��jk/*���&i�]���%��`��h��t�p<2p�PY�	0J+����u�t�$��V���9�]�~~@���T,�MR����p���i���]��Č�<�K�1�R��,{ ˏ����"i����~��K̰��������M Iq�I�wC����,ak��s�P�� �~�	j�qJ�
�l���v���W�O�-�[AN늼�GE�a��m��㈛C��J��w�6^`ɝ�,��|N�]���35A���=w�\6sע�{��n2�΀ Ћ�%���S��)S��K��g�vԈ�n�Rr}-7'z�P�y�m#�}�^m�Vv@�W�և�0��-ɖ6�ƛ@0߾�����^v�z�V`�6T\�z�%�	]8��l��[6���?�p蝫��;����z6��u�]m���G�*��I��FVw?��"椢�c��~�H[)�\Q��ر����r��}�%"��:ǃLt�gj����VL�^�d7������O��;;�LZf)t�:� ��2�!Sd�_.�cfa.'������ �=/���^K��><�஠����r�/���X�j=l,��N�s:I��C�&		�m	V%g�Z�~Y-��Bh��2��ε/+F�Q��D�9C���m!�7�VĂ�[ᄏ�V�"/T[���1�/!����k�x�Vrk>��gQ�/��o�`�k/8{���F^�65_����|�������֦L����х���X��2�J�c������@<C��RgQ�P6
1�Z��0'���$h�k��W�Xi=��\����	���������VeK��+^m�F�����{6�|{Tz|��I�ŵ�
X���j�aē�� K)�xfЮ����'O��n�i߷Сn�d����t[崡�>�ɟ��>`�\E�^��T�hC�v��^o�eC�8=��h~�*�)�����	c�l/�-�����tH=
@����ߵ(��P�/ �0��.r oEqo-Tp�F��E��5g8m���pty+b�ʣ%@5��J�ũ�3R&�9�SR}�7sv�����voV��l��J	��t^6}ޚ!��rD!*5(����Ŋ/���wv��6�W��w��:�[�"!jK��
��*�3�����4isuW]=��
�T��h����hq\D���<�˾�d��2�����g�1]=݉E���4�)�F�	,�"�2��)5y@aH�Wt�J3:�Z��3&p�!g�RJ�����ݨ�*,h�'�������j)C�?�iR:s�t���o�.U.gz
(��<�^���q0p���B)� �Y����t��e�b^�H���e�*вi7�$`P	D_�z\�.V���+i��mS��$C�f箲v5��>��"�%�g��	��ƙL!=.��9�G�`�+w^i�����S~�DR8�~�������G��}���=֑g�e�G$���V>�Y�NV��ec#{���G��͹�T�@L̄�S�h����<����L=W`�ߦ@j�����b������4֓Κ!-A&������"�~JJz6Z���g�x�=�0p}�9��{��g�����-t�C�e��w�II�܆�ԯ4�yG�1���9��f!���¬Q�L~uXUk�਄X����q����,}��\:Y��4�M����-+�W�R���
$� e�7�~���"0P��c�U.6�I�6:�K@���K�t��]u	��](�P\���7�N|Ҍ�^@���� �
��Wb6;6�8���#��:�VX�8ҐjR�7��Uw�31��F"��O�{���I)�� �m��_�Xxҡ*crz��e �l.����y��ڑ�\	g��V� w^!�Pa~-MY��� 7BϞ}(����ثbʁe_������
�����Z>�qDhGq�.W�<>)3�AG)%��-�$�=b��w�CU��&*�>�p� �8�A�3�hp}#����d�XA��1�Z��u�
�l��_��s��C�O��FD�a'��7ߐ�c������X�"r�Ev��2J��-sB�zCD�X�>XZxe�zu�*�
�s���S�א�G#���-�p�������jsUE-�\���%II�*��S��2�>����
W�������>A;��qL��ޕ�����*@hI�o���I�?�n�ukJ{m�g�5h_���)KF�7ا�W��@ԩ/�r�Ίݡ@Q�"�g4��ϑq� ����71-Oa�u��i������O��4U��\M��+�p�p9@	J�4_i������-�_{�����%h�,��G\E�_�?�#k�Ă����d��0����V� �R2���m�Tғ�/�%�#!�DqG�_�"=]&Ͳ��S\��WM?��GP��_�E@�&p�y��{vߑ��@*h��~��#���L�H��@u�����w;�{qw��٣\͢��e��l��)��⏘�ֱ)����';�2m��ጨ�F=��1N�͸"O�-O别U��:��p�U^�{� "�CbɃH1o�;�kv�0�Q����`3�i���OG�~��s�a�򅨍��=���Y�'��:o����V�XA<�4��~�4�.�JN�F�ù�|��G(����\P%�2�D��1��8��b��vINS���݃	 ��֕ː:���.��`�������,����G1��^��	���8A>j�uo��$?�\��<���=M�C��:x��p�p}��oi����1��u��(�ܩ-�XTۑ�}�|:����E�
�>F�����cz�w�zE��.O�VmL���x�,I%�h��0�Q�;��78C�D�g��7��*���U��"�u�;����g>`����(,-@3.AX�=_VYDL�R*nR^~��)�-u2�o4��cݩX���P��*Ј��("I�``	 �K)��x\�=�l��-���N�m��NJ�D�P�'��(/6d^�g��R
]�sL���:��
�x��9~ޒn�E��ut����}u���g��$:VH��ߍ��@�[�%=һN�������4v봎0n��;��i$������<��:*]�]]�SL���K�p~�>)9���,?>Ñɴ�K�C�]1�j́��K%����s�z{s��y��gZ��Cp�x���M�p��'���76���ssi��0���BMtơS��]�ÛS0����~��DG|+�+q[x�Fn�Q�����{�tƚBU`��y��]�1J;�c��)aҍ2�����D��&�1����?�%�G^d=�.d8Y�e����>Y.����CrZc�%�"W�G*_�x"��͜���K��h�e7῁Ai�Ye��mq=�t�����9��(G�I�J�&Y�Κ�D�n���ݞ�����|myH��ְw��䧝[ˬ���=�836��,�镕O��0k�Q�0�Bo_�(C�R�����q��Pr��</�5e�Y��Sq��[-@�;}67�3�1>!a�Wb����ItD��Mڸ�#�ǐ��k�|P:�����o�ۅ=����=1�����W��� iZ-giVd���;x�(�rϡ\�m�t��=���/79��ǟi�0Ƣ@�1(��T�>d�C�����!���B⮄j:����N�٭Ϥ�F�
�i���S'�L�5
Z��U���]�*o�t�hd��H@�U�j?D߶��A�I?#�gIm��*��r���J�P��Z�/��.wH���LM�[*���-��u$Z<�2q���{��b|���*j���G�֦ ����{�`� �F��`Өg:c1�wۺ���z^D�!�R��.���뇸ǻC�<ZQL��x�Rs��p*�'Ћt9a%q�᜹��1Rlm�]���{d+WL�¦l��i7����	�4;^$����9Ԕ_}ST�t�5}��Hx0_4f�D^O:'�Oc�Pd�yyq��rɉ���R��s��?�WX�	����5�)�J.�`�	����'��8�b)0|����gѸ�m�+F��~��kF��%��eZ���Y�T�i�g�C��M�W_���!�Amxq?���@_"X�~��`�	�
��j�� �U�DCa�^+6l`%d	F�C��&-o��xK����]ܤ�kYD�~_)Wi?2�tzW���ҫ��4x��,�+H�0�i�)�!��)s�} {���.Ә.VȵBz����ӯU0�2W}@�HEO��z0���G
�a��X�,E����u�OpBUe>n��tp�>%9�à5y���ԅ�F�����.\�	l��`���Q�b�]� (��<Ыg?��]�v0���11���&�3B�F-0,&� �t���V�8p%<�=���jx�F{��iVp�up{!��G�mlOz�^0^�WE�R�
Hr,�;#�Ҍ�Q���[��|F������,W�{��)X��~hh��������Z`�Z���V(�|5�X	����G���)5�&Ǐ4Ƌ�C:�*���ZZx5h�o���f�X�L�����J ����x��2��u�*�Xt�%��-����H}!=p��NGm��𯯽,��E��k;�����������.JaTƎ�F41_{�'�u��+�/[e%7��F�*���*�T%W�����h���|�P߼'>�0b+����l7�=�q�=t�-��ā�C��G�'E�\��F@nvFB�.�.�bԝ�z0¼��).�`��Q�@��o����6�%A���⤣�^է��6J�k/n�eΌ�(<�Bi&�uc1!�)k���-�$�
q��S���tޑNY�e����3�g�ʏ
m>�Ȍp�Rw�������.&�&�Cu���{8��B@�F��h����B�9|r�D�Z%-�(�G�G��"$�aXa��rA��ں��V��Ĺp2z�8>�(����Xam��E$E+ga�����fs$����x"���v�7e�ƸTX��x�)Jz/R�}H���҇$�9گ��^Cr��Ӳ6��ę����sv������oXLdV=��,fg�ek���h`�@�db����/��
�ҍ��+f5�L��<}�v�@�O�z�!Z2��XCm����Q�����������X �GL�,f��$`��0�E�����nZ��X��K��G��Թ�Bg]a�Q~�7'���t&*��~e4�7���ih��o�1��
��jP2��Oi�mfA���(�J@>xxi�n��P���^�}���I�"Fx'�c�R~2vd�їl ՊF��$�ѩk���p����?��p�i�WwH�'��^̨�|��^��PM��T��)��b�M��.J�I� �Tz1�ѕnou���d����"B��R���ݸ��Y-�	K��P�
�#�f��U/VZ��ug����A�xH��5�!3����ܤ��L8"�v� �����tl�����D[�E�Ur[
]� @y�跳���=��U���\�/�u�M�O6�*�FMLVv/(��(��(uwJ���%y��	��(�]�I(����No�ri)�,gl^z[�t�lۼф�g�P6.�aa�^��@N�F������S��6�{o#�xYM��ҁ��jB��)��^Ӣ9c/a:� K	. ,��,4��;
����Q�R�
�Wi}`��T��%`���KlN��C
;}u�U���5�n�v��W�Z��:yE��E�-}� �����4m��ɐT�*�� ]�1J⮶��kL�7L9�
�b�0�9�eUK
"J*2��2��6�8e�Z�T�Sw��K);K��@��x]�SJ���5�c����*�መ���N����U���7J�Z}3���#Y�=��j@���Vp_���+L�������L{5�"ד/��g�����Y��yd���E����Ge�m1�p$�+�Et@]'W�*ۚ|�����j3����7wGp�;�>�=�'x;yQ���|oG����`2B�8������f�[��q&��d�vC^���Y?�F���=	A�T��A4�g�mĪ�q1�*������-��r1�)�6j���.d�~��t�xƆ�/���3|�@�4�e�z^z�����	�J�cG<��=�Kw������M�_��/��%-8\_��oUH�d�0=����$�������Y�w���/���B�gz�uS\c�9��z�k�-�`UnO;���j�+�y Z��Y�$���y~�Df��<��]u��e�B�i�<��I�z{��Pi���@���E�Q�ф0�Nw=G�G:V:�0���ؔ8�J&q�熅�4@�צ-��d�$p��y�}�3�;:�W�Bc���2!�E.�A�Lz4�C�����p';�`�Ҹ5��1D��6��F�im� ��Ӯz&���{�_?xP�B:�S9D)n~�
 ��pK�^rY5})��c�-y���5��p6L����{H(�����S��0QN&W��{�~��i��n�����kNi�9��Ѽ�)��y4*	nʝ�iL��ZV�2���5"(���=M��'h�:bkT��mN�o��>J"�q�;����L��^˺Kt*Vǩ�p�w��#U�
�{��a�U����e���]�A�������<��D��%�& ��Q�*Ե�	�7�w6EU��f�u;�5U6)��b*�w�ƑX���{-�hj���v�=0l��i[YF&qX�2)�F�v�uU�YL�����`2���y?�YW�}��]��N�tr����D�qO�X���S&�s����U�}*S�ᳯD�6�+��SSѼP��d���!���Tz�t���먼v��%̎�h{�Wl;3f)�2ٙ����ī��o���(k�M	>�<�6��Ȃ��{+�
OȺH
b���Nw`��D�Aq�o�^�b�+�� �|_|kuB�Ү�����Ш��������*,�d5���L��i�� �H�dR��C��	�T0�Wf,��j�x�e����^�,",Z{��_ӽ���Ab�&W�a��4=��Y,��3�2��h��9��N��%�ٟr�S
I�a��Ӳ2#i��=�+�Z.�["��&d�tr�S7��v�*uJ���))Jj��䍈ͥ�VH���E]L�L��UAR��G�8�h��4�s
F/�{��֩9��9�c�Y3" �]�_0�^�]:yߏ�+�$h�x�<�i��r�˿��La�Q�{۞L��6����HsE�RKk�!��ZZE�wjf��Mqc��9���6¹�R��<X�a�s���٩jL����O?�1t���3��{d��bX+��R�OV+�!��Y������N,������_�-@"����ȾX�f��sFV��00A�6�S6�N��˘s&.�3`���02�˕6?�4��uMTWƩw*"۳-#!_jP�-#��.��7ʟ���OB�9�>���D��|�Y2��Pw3��&�<J�n�%�&�ڧ�O���Q������l=��`���d���.;�&$)lk�U63�9�)��#��褂��)��.-���;}+�7��B�45��������eA���������)&�����Y�]*6��+GZ�gp��	ӹ����m��d%2׭��,���R�I w`-f�����F���~Zv�������D��],NE����}�s瘾(*������L]�x|sw�&P����8a�F���<~!�(~���!�YS��J<�L�r۽T����M~��a|"{��i���'�e_q��%I��c���%�ѹ�p�h��ڼ����
��������E��g�4b�/�Zħ��,�,M�� �
sEn�fZ߆��D�{��`(r�h%��R�d�{��������Y�r��-P8��Ӄ�U�%��T���Dh�������Q�k<鿐�v�P��"X���	ۉ��K��>-�0^�*�=D��f� �?��>���=��9���������X�R��D`�P���H�����g,:¿�y����N]����!�PC�,��M�bQT]��Ÿ��rԺ*u�N4�So��_�j҂�ш9�8�F>"ܟw�>sh�9@c&�������a��̡� 
�����#��9��w�*<)�����"��q��veI5�5��_{1,Q�ǈ�u�vX���z!�e7��T����I>?��o��;&:Q֦f�Z �Q�Y֏�W�*�W�t4����3�`R�t���9}�&����:������O��D3$��f��o�,�&��ҡs�F� ��>�T�
W�R�O�{��3�)�a'Jl�ٸ�_^��T�q�Ə�5�������^��Z�V�y#�ZK7/��+��W\;���
JM�����`�3�u�������͸h�qA���>�7�J���r�,x/!��m�ҧ5��o#
�hy�t@Ab���p,��7�x�)J�R]B:��=Mo8��i!�o��cw��e���:���8��A��2�B?�h���q��lM��ch�g�w�*~�T�E���u�5YG���9��؏r����x=\�3B4O�՝GV����^�;]rÙ���+�Y`t���C��cς��b|"+@�$�q���0?�������
M���:��[1X茰��\��BK�r�z+�($<�;*뵖�_Y��۹xU����mK�z}��[t��R@�'�2z@U�0���a Q��^M���'cC5�� ��M[O����
ѫ`/������	º��\����]#޳{I�!e��FIf����/8��jwԒ��cjetF����jI�i-bC
����Yq�� �͙_���e��<��p'N���x?�ڂS<��g
�z�����Pxb�|z�nI��2���1���-f:^)z���NE�I�����ǱY�}��?��<�{��Μhi��ؘÊ��cq������<�Fo%�y6j�a#���GvS�n&g�<dHs����8�s�SXh>��!�c��&b��8�+q D]��fa\`�&V��w=6�=�h	�����3�R�M���bȕ����	�$��p���l:����D�E�V��sp���pb���4P��!K��;3��&6%K�l׳�[l�P�jg�O=���n7�8������wz��jx�-p 9ݒ1�l|eη�5|!��u��U�����4�R�C2<h���J+s_&ɩI���O,�Q�ӧ�Gk@^��D���gﭮ7D�<�IfF��%���ܪ������p�刨�޼o�jԺ��ZάQ )����I!d�Z6�����(Y���i����rm��}�G�#U&���FŹ�Jؓ&�����0�{I7���8A���K�#��e],
 �m�Qv��~<�˓37�{�$����;���$[��?l�`���8�G�������e�;X�ԱGC*`g�t��GMa��g"�B�hc0��j �y�o}��D�iZ��D�HG����ٙ.��h�.�7}�Y��}��D�����l`�PN@���T�W��l�.�qy�o|���Y?F7���NGZ�?�Uܖ���8V�p7�.O܋i-҂[Ju�-�Ƥ��̑أj�zOJ�g�S��4F?Q������w�@�x�v��t�G�9<��B����g��l �h*�YY�S+� C�������`Η�\#Uj-C��XV�%B���w�Cs�O�v�OpR��L���S�p��L��{�
2��c􋘩�A��#�2�#��=�~��x"�Z��I�7�A�$R�����a��q�W�!�w�z��՗o�@��(]:Eg���j���t����jl�U���`X�Y�9R��5�|��J�s�H�����"����Ֆ�x��k	`*�&Pޒخ�q����X6�u�@}f�):�oEpPl~XW%�M�zCxW�Y���}dq���oȺ�Bn.*��%���_gp�i��N���%#���E�y`&ZQI3��L�S@�8K�#�[��Y&5�]v<.7]�
P<�����m�{�Nz� �N	���1&��Y&}Q+��S@-���I�Qyp}�w:����gE
��������dS_��	�vEqE3�3ܭ��n�!������Zc���58�L|fL����2������T����c��.+��=@�� v�,�y:X��F�S����<���ۭ�u�
h����S@^�n�nGxS�ή��4�Ǿ��({ƼH<o����Ʈ�#�o�i��ܵ�Wﵤ���%�~�fg���g�?<�3�H�L�"����G�5f�^�
�e����A��J��������z����wB���	M5A��5"E��h�u������,f�+:�+o����ы�������u?���J�Y]o���������Jz���|�U��%$���q�ؽ�H�g�\�	���׻�"�c_mO�}Y��)%��J�b xn��{U�`��'yt�����<��v��>+�7/M�����M�zٔDO�n?�]�h��[���JVq,۰\Y��4;yK֔5���p�'�EE����$v�I.TL:%`�[�l����p��=��uQ��=^p���3��_%.1��� �Ώ����<9�5�R�-�A����0W�9�ŻM�ʢ{�k%/� �:�Լ�Y;�t~��,�v����I� *2=��(u�8g�S�
X����-,�P�UB�6߇�#��S���R�BG��9�}��%ϩ2�2"X��3+�7&����g�ƣD��p��X�Xk�H=��N�����7Ns��H���:/�v�J�Z�)����&�t�b��-�(��X��"U�S���_���̙?�0 GLUnK��.6{�%⽎)%���_V�� ���k��=�vQ�����{����[.������!���e�"+8�h��F�����Y^]B�(I�,���r���	0��վ�Le	�߉*����f405w1�a�a�3"*^�<d�fso
2���dGa4T��C�v1���d�f�v%!�K����:;oѭRU똃Zqld�b�8������Z�+�E)��K+�87���s�'4�8t��c���"��w�
H]ߪ�?	�ˬ�vM8��;z1h�\^z�2�S�n
p�/�_=��8�	���Ϳ��{P�W��Vv����?[d-'K.u8qY7��r��r��:`
*$\Q�e�#�(�����Q���mK�s�M�1�4ҝ��lb2
1c��������A8 �]kl����Jm�����J=�=��3)�%���ݛ����������ng�j80�mLXAe�S�����Ũ�������|����N����g�J⏕�����ϵ]�,�"�\At��.�z���o���P���Ec�te�����ʌ��t(��g��I��C�g�s/g��y�q�=����P��ւx�E0��M�����&nhJ�dA7*?�����1	�z���#Zv{DAi��?���������J��#m�[N0��#�aI4�a��-�Y��8RV�+~�	'�^QR��V4l�Q�d���Χ��X���z��3��6=w�&�7������npU�f�Y�-����0_�#�� ��j�F-��3Q��b����s̜O#�z��`���OA!���y�n����'��?1����U�j�M�I^���W�L#+�Q�)N��
��)�.�̜��nmD��n��>����U�	F�S�-��9>�s����s]ڧa�(-;g�G6�(�Zu#���W�q'�^􈵟�ހ�eߔȴR1�d0N���pb�>�%1��b���5��"����}�ڐN�'�\9n���V`��+&7�cy����1�L�}���$e�D*������q.�w$��������Xx������?��kE�f�gc�r������M���i���٣�-MܞR�GZ��4X>��������_�X������M���lv�\.Օ�9��	U}�p�q��>DCM���b���D�߷�X�펱r������/u 1��yk��t�q�� r~�0����&,�k�T�A!Z�+��� ���ԁVAQ���P٪ 0.�rT�d�Ԟ�IN����u
[��wZ[H�L~M���.�`˻�Ԃ�!��+�G�J�V.����i�|�{)�R7T[&��L@s����pH�A}���Ċ!�fђneP����d�dj�Z���d�ɷV E�xvpO4��D	��/��@�1E�+�Z]o�o��sPu��E��xY����e�������k>��d�����R'UX�	�Ǚ�oB.�c�^+��p�)��\T�$^�h��|A�&���VN��u��62�b����b*ĉup��& ���K'�6rD�q��o!�hX!6��e� Q�h�A�5�N���9��$�8{��w/MBg1�n���\ݺ+a='�Qx�\���ϳq��*Q9K���Ǟ��6P�iɧ�r��Zʓ�;��3�l1T��K�PF�:�B'N?^�p?:;�x��0!}B@��Y0��z��՗>Prk�=ii�@ Z����S��������iQL�Q�ǣ�K�[�6o�u��p�C`�\~����Cy��F+J��v�{a�}�G�,	��-�aᗞW	]N*b�2���ˁ���g��6��/�ˈ	�&��)������۸�h��F��FZ�Z7__�T�o註��'����AX��W!��&����9y`k�������Ț��(��z�zA��򿈋�\jKq	}�Ux��ٟ��Rq�<P�<�-�BS��>p7(�b�7r\\�G���������PAk���}��_�b��낅��ԏ	y����#��>���F�2w������2�:EdZ}�7��P�����iNםLã`s��s��]x�������TZ��K�>�����j４C�b/�=]�	��ԏ�Lp�W�u�r�B��հj�b0���a��;*NJ�*m��F��