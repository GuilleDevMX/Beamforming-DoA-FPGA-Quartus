��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C��(b�g L�N�W/u�b|���@Aw�_��5����w��&�T�`x��i�>+�_^�u����V��0�d]���v2�/O��iV��'&����%D"[���1�����4��b���jEv�w2��&�q�%�fΚ��8�n��_�fצS�
D�aA��SRÂ��߈]h��`5K�����:�6!]�9���6�e�?���Vu�N
wش��Q��G��N��8�E�%z@L��"ؑ9�"�17�%��(������?���}��[��81�)������
������(�mv���jVK�`�O^M	�+:�I����z�x�1/���È���?�(���с�fFƾ���Y��D{��R���'`�Z�ŋA���(M��+���9�%=˪0�7�5��\���Y�`�L�
���A�x�J5��1W��o����
� ��J*&��|�L7W��uç��B�(���Bؼl̴���q~��a��K"����b���]xCm���W'(��3��6�&�!��r/�*������r�����h.Dû��52Հ��˳;��B�c.�a�����;;���}�F{��oP:���Է3\x\�djUr�~��:�� �J�� ɇ�.�'����^���m�A�@a���<����u�2�j�5���h15�Ϥ�xl����8B�]p�҉�U[��Q�c���?���SK�xG@L��S�ڿ���kw�(��!�S�"g�׀�߶kG�f��Θx2��a3'�(�6�-ֳ��n�㸆���Evo��і�UNL���^�ǁy�/8;op�E�ǩ�40�J�2%�C��r� Hd�׃���)�y�,�Q�]��"�p��K��.�69瓉�Ǳ����}+z��RÚ����H3�1�{_��swE��yP3�kZX��ڙo=�7��(/8���Z�cq�;�� ���}�	A��Vö9�L��n��!���"y�.�XK蚰����5�|�-��A/�Y�ʚ$�I�E�|�L4B��,'Ȱ�c���Y
�>�B����Yq�y�2�J�[�|[{!��f̸HM�E�R2��_WJ���<�g~˘�v<�{��2�*W+�_Pc�J�2��� /� �v! ;������"�t���Z��ۆ]��J��3�	�0n�`��hx��PC�<��؅��[M� E�e�d��'_@�m����5��
���11A�V�o��_?�?oj�?W��� ����D�y8�[�84<�T�/�x8Ɏ���ψ���rs���ZE3g"g�{��l7���k�g5Vmi(J:k{�$ؽ�|".�K#��#�����b�sJ^�����T\����T.�cI�2��,FPc�ݲGZ���&���&�юӒL�x���}�w
.��f�xL�d\}2�{D�RC)��ƇL�S�.>8*e̞�C��43/إ��§W��k�3ӫ1����P2�SqBe���0�<ݟ�7���t������FV�?�3�A��Ty7����4���p�o�԰� ��N��!XJ�^>���g�������W��+�u�ȃK%K�	3���#:++�sf��N�J����\���˚���G"�h����`Pw$$�ř%־N:�ĂU�_;��#M�d�z2�K�ԺoQs�=B���@�{n��]Z�o��7�:}mBh�(���*@&�,(��1��{��F��v��ia}����>%�"C�x+e7�C�ڍ�0!s/$�M�Ce�����g:��t��>~ +�R��M�O�uTKׄ�P�P���W�����"�nṾ�(٥G;F�/��Z�-�0�y�a1t�g�@M�y�.���e�J�j�O���*��o��6�a��l�A(V���x���ɵ�
:�9U�a�Rho�?��-��oI"�͵��W�w���a����釆��n��+]�2eWq�������co�!˟7��&7�ʑ,�A�C�SM�2�dS8�Z!n��+��!C~��`.�az.c����3H��^�)���6k�5����f��V�����̝�j tS�=�V*��Ô1c�)c�h���#��b܆��%�u�~Y�4� ���Ե!���䵏��>�a{bpU8�z���j�Q�L���l7[��O�en�±.�1�>h���gsjz	�8D�;O�,�uS+�7���#�WD�����]j�t������߳g1�>Y �AN���s�.�"@+!� Ɠ	$�-����x�?!��C��)���wd�j
X(���R�*E��}���^�Y{�br��ȗ�˂��*cDg/�+��Ca�S�鹬��"TgS``��-�v!��j�	�?��$齴d�}�$�=���$(�~7؀��c�N�����g���
�"x����ң������t�
H��TQ�ߵg\k�	����ێ.�Q����+�1^�?F��O^�N�:� J_�'����{*
�;}�Whc��y!]�\.Rլ�s�y,P2�5����Ҹ�7�u^�<*��nކ���11���W�*���Z���c��IJ�c��i|5��_�p�Xī��x�6D̸sB�7�pcb=ڈJ<--���;\�f�Ө�i���8H�~��?2�7̘�yk�(n��_��I`=��i�l���F!n�lN):����N;���W�j��K�Ij{���Ԟ�`�^��gk�$��i��i| ����l�=l���B*8ێR���󤫭ݻ�Iԩ`�S3�!�K��%*A����ĺ����������ˏ"8��*5��L^���1��@R��Ё�f�o��j�/��p��y6c�tD��}]�j��lz�_�7��<�:���Wn����}NZt^ǅkCN୰���7<���]<�M�A?� a�trf�Į�$�{{�7��`��X ��tL���K���0�઺34�Ng��_d��@<@;��������r�旣�	�jd����slf�(8 �akwc0�� 0G)�I�M��5��2�m�u�'g��~<��b���LTp-JfZ%��/�|�o��w�<��~��lZ�ϻ� �Y�����ERXw��4��a��Sf=2���y�����ɓ�\<���T$g����k��٦s���l��%(h�4��[�brD�+>z�b�1
T��V�+5,��(��	�ĵ��
�Г�mwZ��&�W!^429=O�l<uzI�Q�s]cr�K"���C��(u<4.�����zp��ݡ��Ǫ@�9�K�lɷ*V�M�T��٥{��*χ��z8g�O�a��T�jcX��52�}ʌ|t�����7�(���a|ǿ�}�[�Yk�z�%�.-rᰆ�ݏW(��l��C������'A����2�)t?{�i�h�X��K�#t��	�Ж������v�]�� ��H�?
����)�[��V#�����O��$���jm�X���Ě�*�ޅ�31�q/��Z��v%ڮ������l�b��]F��hDv!�Z��Tty�r��#|K-6�SI�J@�m�V�uӖ���VE���[��!,�c{���0�մ��*�������P�8�22/������վH%=���e"{��R#����N��;��aUb��T�o���*�^��/,*J�_F5�Ȍ+?8��#�R�KW�	h3���7梵�ayM)�o��^��Ȁ��Xz�z�;���v����j̠cIק�������S*�/q�^q*Ч6Rc�r�A�z�tC�[��*�
��T�����b�=�pl����&�u�F�j�薻?�ݒGy��ӢO���\\K|8�:4)�O��.D�쎈������@���IjVق���7� ���/,���9	�}_�m��ZW��hw`R�oO��b�����pݓ�3�����"��g���N���GI>E�j�L���$�}��TN$�GG�D�D��q5�YFTB��k�� %}�^�:{�a�� ��D�)��O}L9=���Ѕ��)�j�K��7��S�l%'����W����x���	�Ng����_�_�Y�t���ֶ��\��W��\��h� vT�����'�;�U�#���j�V>�Ѥ�l�c��,��w�6�b95��_�
s�b?R���E�������<#�IO��TW����ވJ�@;��9��{�8�Rؠ-��4��aֵ���S����Z.`��[*���n��LD�]*�⦄ʮ�41��D4Ќ/�W�h��,t������q��\G l��E/�x�z�:16��Mbۑ%�G�
�{@3���������Ï'�������QG^<�� �:Ma�Ȓ��!�0�e7=;O�{�����w���8i�[��<e�x&�X�kn�F�o����M�Y�)��-���汗#�2ӿ��P�D��a"�P� 0�E)N�O��>(�y�3�^��8)P�!Ad�j�V���Ԩ�x#K�}cՔ�.#V���R�����a
��C��n̟����QT��_�oHp^��q.~]�~�ǵd��`?h��0���U�"��/���O7��uB�G��?.Q�`�xTɁ9P�6)~�L�a� K���Pc�}jo>��YC���|g�� ܱ�C�ٯ5�G���5�(�} 7l�\	pR�m;4�!S��7� �C>us^�֑݋( Y���{�6�/ _�����`���vGda33D���7�RɥŬ]��u�fE��׳�""��t5��i#�G�����XdS"z8�$�u��Hj\�mJ@l�0z跔?�)U�`{>���VB������6��ߵB��ufa�f�^4�����\�ī���E�Aе=u�:���oUd�Gw�T}�㊯l��J@���Ɇ�p�C������F\i52�
x
P���~73={�W��]���L�hf}ݶ�A��褦<� �_l� �����n_梂�K��$������.�a���i�l �'�y�^�Թ�}�r�ƿEv���>����r�P�>A}� |�6�x������dU�S7�v�k����d��!��6������FآU�!cԢ�K\���(jy�=3a�������������I���!�c�bs�A
{$�_�`��jhz����!F}�g5��.^ N���:/v�g�Ԩj�rK��1dԳ��h"�E�@@�xEB!�kͿ�ӻ	*�q�A����v��׮��:��䚯t#�����5���}j�ߐ'ɵt�h�l	�v�,��X��g���x��	��i�����]_t��L#%F|��֒`�������V��?�k(h�cRO6V�få�29>�x|��2	�:�E�V%(�׬��I=�O�[n=9��ui��;s�y^�z�d{W3S��̑�E�j���m�����㨏꾭��V	U��y��5�̿wy!U�vQ�쎛2�8�hΚ�%`�v�۸8��ľAedz���M`W`�M�f!]S�O����1�f��Bg �$�1mK�._>��j�ǻ�_�����ӮQ5рx��^�+��-��f�!���?�f	����i��D��K�l��u�[���Xv�l.�֐FM���<6��d�q�I9���8&���U��! �\O�x`��9�xYj?9m
\�X�γ[�