
module serial_com (
	clk_clk,
	reset_reset_n,
	rs232_0_UART_RXD,
	rs232_0_UART_TXD);	

	input		clk_clk;
	input		reset_reset_n;
	input		rs232_0_UART_RXD;
	output		rs232_0_UART_TXD;
endmodule
