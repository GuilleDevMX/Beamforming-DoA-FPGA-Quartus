��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#�=b}��u5P��>�� Vߺ�D���� k�gU�n�P���ِ�+ѱ�{e��^���g�@���KrKӾ_z
�^4�z;O��T�Q������d`�ں�Т{���8p�Kt,Z߷�����'�NN�?$�jXC��Qt���;����HY�L@ry0���&|�>�x�ڑ���#
XA��#MI��ك��djk̢�L!�g|���<F�^��l�3�1���-t8G��πG�,�r�e��a��?��>9����권A��;bE��X)gS��VNGP'�5���wn�[q-��jla�Y���H�T��c$Z�d&d+�q���>9���m� ,ӄ�&�X"�/y[�w�Y���b0�	fJg��}CW�����;���v=��4$[~O��̏���$~��z3G�ۮ�,���;2� �O�I?���$�YTY�B�zex����TEQ�5M��Z�=KYX��'�++Õf�[HZi�����������f���X�V�m�p�a4��!�Q����M�	��9��E�c�>Jt��r�ͩ��<���.�Dw�Q4��i%��N�P:6�0I]�9��I����m ?42 �C��+:̉���KO�hù��ƶ���Ѧ��ϼ��n��V|�zp����mG�wȘ&�\�|r;�!n�~��H𒼄�井櫩,�� ��OX��vs^:���9�ܜ�2>�_,{g��oUH���ɧ�xJ7��你C�j�v#b�"��3{g,-�xT� ϧ�jC����O��X\_��>2������
�S5�j�5����q�J�UpJ~�ԣ��#:%|����/��V��#��7	�q.�'۟�6���`YW)@xBt8O�u����}/���b�7��cx�A*�M$�7�l��~H*U�]i�a�/[�b��3��@[�/O��E���D����d�{`�:�!?�;(���rK��(L;��S#Ps��]�8P���U��Β�`�y�7�R�_�"�|���h�oRG�C��{|�zl��5��Ou8q1�{Y"�ko/�@�Q��C<fo����?�	��h&��1Dg��c��ɒd3^�/��";�8 �m�K�rM1*kc��$"p��T�����n��.u�I
�6�=�����Pn���?���#�_�P6�H��v�P��!pP�j$O��8j/��/m3p�2�@tu|�iGq�prQ6�x[���C���eR8��,*N��(�d���_����f�=��)	���5��`�g}�*:pugf��g|�؈7tP
,;��c z-��׽{(�.2	3F�cVy�i�=���qXbP��iOg-�Q��0h�G�*�E�-�Z�UWo���4Q�[��E;۳�A�I�Nc�����鋦@P�1����1�;&����YP�F�p>Ġ��2gEr�O�:��%�g>ځ��T�!�u�U(��j+���\|�f�ː��>������6̒�P�+N�wHU�
�M�e��}|�l_܈=��rm	���7����1�~r&������0T�+µJk�V�#<���u���x��c3��5�bU��y�27�{BIAG��yo��wާJ��ywj�j$w��ؿ9<��� �r��
j�F�]2�"hEZ��ݹ�O��C� ������)l�[}\Y��P�Y6��t���Z;�^�7���f���b)�%��o�1A��s`����7�Ej��K-z_.w�wS�F�݆j�V��EN��F�/�ea^��w����|m��'ܵ��Yj(��8~�*O�gȵ��n�!���'��PY1�s��k������d��fO�w���fz_f�����_r�����7��I�(���%U�� ����᏶�*�t���j�p8vU��l!�7T�b��nA�ůgN�R�kT��1(�ٜc���s���\��-��H0n����z�7-���x��#]۲}5��us����'��eZ�R��-Xg�=����������?2u�ܘΆ�t¶�e:�����M��j�$�P��S=̘��q�<.��6,J,a&WH�z��S�ja�T�gdw,�M�d��D�PJS}a�8gŪC}wz�N����q�`�^@��P�q�\I���j��\S0����rқ��U����-��DIW,y��'=�Fnz)]�7^wR?�M��6�	��yJ��l��~B�	�oFʤ���Ո����\	�]�r�s�c�
��&���gu+퀶�b�i^LO�H�h���s�?�����g���*A�T=e��Z%�N����q��b�r�,:�xSʷ��	@S�Ģ����%�GE�+�H&��R�?['/qRt�s[l`�7k(`
�4����8ӯO"�ZZQ���]݊y�)���/)�uekUx���cڥ_�KCT�5�(Z[Y7 Q'Y9qʩ�e(C���5*h���.n�x�J�sأ�>bѠ�o��74ҋyQ��� �5ς�����0�3�xG��3%P|��&"��А��A?GV3t��ҩe�W�# ۜck*�W��Kڦ�7���"H���-�,Ci��X�x�_�M��'�~-���S��"68q������% JƂT�M�<��&;dً5DKn��~���&�.�0 ˅ϻ�~� ����&R��^;�=�W܋Ɵb�L�#��D�֯#�-5�h��J� fXӃ���{��7ϐ�_�U�U4!
����m�0<�U?�}�G�\#|�0Q@Uٿ��a�O/ؿ����?_'^,p�~7��X�x��n�9��\b�mOg bdfY�R\��W���ҁ�$[��f��d����p�	��ʪ˧���Ҕ�,�'Z��ߖBa�x1�)�#�ҵ��e�#o��J�S�s�<�0��ڊ+zD^J�Vշ���.9[��?z<ۺ����(^�+�;����"��r�ҿ�m�N�l�N�gA�*���Y�e���WV���k����οcW���,�����J�?�`��(��������NuA�fB̂��uW0u�L��s4���i21��Ljl�i�eX�X�D ��؜Q��>�Q ̯ ̗����y�/Y����:�+�s�2��A�R�ܢ��v(MRA�	A�<)���~N�:Ӻ��J�����ӂĝqR�d�S�g�t,޽�B�bɪ�H�LUrm�{'�Wʜ$�c���\��1�/m
�F"�\N�	Wv�I'Ϡ�%ڂMģW#V����ʸ��*	��z /0Y.��o?у�D�@�6��yK��fp����y�JQ�9�Q�	�0�f�����v��Lq׵�|lq�H/�3��ˌ_����/���+��l�ߺ�ݙ�H0�E�ѫ5��x}�];QY	�&�~��/;����ۚ�õ�>��ÚfP_M%q,�\\��,5ϑ�.V�:V�����6 �,b�{�����#w�\��5P%nܚ�󔑤�����cw��Z>����rt���Z�p���Ǣ�}�;�������`C��ӝ=mFc��!"�a��]h�I��{���R��S}�G�s������J�� ����������/�a�B�a�'j^�T�q='����ɰc���L��t9@	
>ʵ��v�p�Ybs~Gk̠#��m�n�=��)�h�7%FF�F�8��2jl�+���M����ˍ?�T�L`B��x~�]�n���F�k��c�����-Z��� *��;��9R {��)T���*M�;_aH����JBj�,Q�J4�p�bک���� �n����x
���L�,z܉�8,��>� �������Bت���q����ջs �?�(��v:�\�ｧ�	�;d �(?<�XA��@7���������:�s�����������Xw��|ԦQ�>����������@�t ���y
�r`!/O���l>?�ͭ�}��o#��O��N3���6:""�����!:�ٛ� �fpq�]�����8IS)8|۞���.�zH���`6_�Zj���;f�Ev�L>��1��t���r��(�Ҁ�ODj�Ti��,�Pck�{"d5����Z*�/�Э�1�b]�xP���)�	ݹQ�S�Y�ڽW.
�2�c��r-��܄ ���YJ��CQ�;������(Q�ðET���:���Qk���yk}eV�@2@J�K�MEu�ߢ�@��,�H1�ߜ�)ބ=N�(�ƭ��1�aA�Ь����>I(n�� �9{����(�>x�#^p�ID��Pvtʹ�<�ԑm�FW��T 'zQ
_���)y���z[����ΠG���Wv���r���h�m囆�Y��+�"�<�����W������G�.���7=��0O�� Km�e���E;��o����m���e�3�͔�w�G=�ٹ�)$)}k��Ɛ�)���&��?�so�Ϯ�w�Ku���^���c�l���\�̬��-}����i��@�u��;�7@)�ƕmx�{F���D���JD�1?>@_ \ ��0���%��8W�`�2.���T3�%}�O�3�߃����7�<d����?��-i�+�;2�����Z#�rmS�<�5�߀�d����oY0^�.���C���ig����Ѭ�~���)�{�h!���\��s&���Ϛ�g3Z�$�X�]U�k������ʍ5�G(���[��e��QO��4�_����Đ@�$��2��֪�2��9{�yEO�$�I�QU�?�Q�^5.��~a����z#�+������	I���ȶ����G�pnm��
�'�`���G9�(�0�$y�9۬������HnW}�v�T��QU�)T84�j�߆�����Ud,�b�Ȓ?�
�q/Dɉ��w�O��I����(��� �$-������r�T8�x~U�>��c�_#E�=Ӻ������-Q)��Ո4"���H^��f�]B��{�n��O�z�����%���xl�-�[U3�J�֡��u0�;�ҳ�.��WO܀d��I��͑�Riy���"�]H��!��¡r뛣������&w{xvU�~����놩]�*��[�ߌr<�Œ�E����cE��City�^݉'�{)��&����2F6}3t,MY�v��d���u�j��"Wn��2ka�_މ!n~�<=N&��y"es6��cZ��G^Ue�t�遃����*�⦲"4�P�'\h	⪄�tYRW�T�ȍ�{a]���_��ѵ�u�$���um/��QE�M"��C�ɘ��"B^ �h�S�ԖaYo^ LR����v��0P�d"dNޱ�h��X �/���F�1�gq	���9*,5h���	y��ƙ!3#�G�n�Y�=�}��G\>�K퉴��v���Ѕ�ts�5�����qI
�	��ி���d��9�]5~�[BM2Y���n��[8o�=vb��ۂ���n����fs'�]���*ޡ��\�]&*^��b�� ��ţ^ˁ�?�X�	����Ȉ^3��%h�xl�=�w
tm!�y� NƧD�t�]�۾�BE�:W�c�#���E��M�z;V)"8�N���Fk���#�1Ƞ�(E�v%�m�H-#Y���Ϝ���<$Ձ_�O�J���dm�咂�r3�5!v���h� wʒ������$����쫙x�1�6���H�|�笱x������,��� �|�r���F�l8�Qw��ΨA�@:���D��u@��~��r����Z�y��V��i˺���㭷�({rt�`5��7,z���0g9E>����� �F��Yܻ��� mu G6�\q�ͅG��v�N-1�^��81%�'��b|byMԀI�ƍ.����-�~�}�1N�����B�钏+B6�cl�W�W|q S��f��6go�*H]����g�`}����X�0���jY"�a��@��_?�{e�W4�EQ��}A��\��/�akv�&oHf����#6*X�ݲUSR�Be10jd�L�	ۅ��$N>�U����%�1�OaF�vN ��Wby��sf�'�>�y�x�}x7-B(��`��M���g/{6/�9r.�'��5��6o���zC��'��$F�V.��D����H�^]$T������+y0O����C�-J�T��8���6k�� ̷�6f$�L����&�ױ�E�q����r�o�� GjM�]�.��2�����R�q̉��72͆1��ԙ̋�1d*Q'� !�.����Q�/[%��3\	��-���e ��W�������.��A�4웕��k�>����p#�y�s+&ڀ�>���`�e�����o{��� ����q�NQ�^���v�y?0۹��/�=U*��?Ep��3R�]{�ˈ��L��.�n��a�bȲ~پ9P5P�a
y�]/��31��n�S����?�v3�Al���a�SH���=�2�=�3܄�=�ݒ��