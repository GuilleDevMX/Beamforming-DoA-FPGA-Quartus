��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��|r�j��rx�AQ�&�H��F�q�(ޏ�a�K�fv�d������������4-1��vɣ�e:PSo��+�fW-�O �0J�&AY�`�N�����B��w��o{\y[!-�ZC9���~��{��|�G���5�[iN�Mg_��sL
�H�����Cٞ\b+�`P����>��Sߧ��6�?<;)b��d��ht,JT�����5���#�C���+>�����Q�?l��#��%�a'��YTo��q�%#&;��; ��ZN^E��`y��Q�R��F3��Ma<�6&g�ɹ�Ɍ��A>����k��Ҩ����`S����`/�Y��ik�$4�-r[+�\0��۴�a�6�l;���fd���p�FlC:1��2�V��AdO��7N��1��0S�[�Hon�E��k�7���������o"�T��ޔ����ӷI�y��^��(�'�)&���8��<�e-B�
�
�Ė��p��;��ux����.���TE�͂�$B��x@>���xN(ց�p,8��b$��Q9yEw�<��E���A��K��(��������D�r~ˆ�wv ���=��pL���뤩I��"�K���6�Y��f�y��v?�9�ڮ�Q*5�8-T=��0qU:�U�+.x�dRL=�$�v<���3���.zr�KN5wCÐ���bNuU4��:���=���A���.���8�.5}ƪ���&"��!��ͷG.�t�p`Wt�@�W"6,+jSVP`hg���|~t���!�XM ��YR��?�ޡ��%�s*��K}�����6�I�7�hFb���L!r(XWkǍ\��<[z8��:�Ѻ2h���k���釯��������4�!7 H����Gc�\�==����O��*;����MfH�Ę(g9D�'�qK&7�������"��T�p�m��C�x��M�iR�������ӌ��ev�쀯GM�n����D�X���q�*�)���N�>N\��KM i����qt ������A����ߒSzW��;����6�� 3?�x	���,ȁ8�b1
C��8��Y\��2���QT���Cgjt' ҝ⽫���H�~�VliB��H'�!�9aR�}Vʯ�z��hMrX4���Ϭ\X6�HK��ˡ�, �+����{l=�4�
6��}�0B+�EAsv�|���Q"���鷳��`e�0��)�W��%�gʭI@���Y]�,!��N�[}�;FH��S���eJY �f�n�[d���n}n.o�<���hB';zϸ���Y)�Z<��������8���J�@����?R����73W���zV�5O�&8���,zwbk���) �^���6�ߤ��<~rn_i��sI�����rJ��v� �4���3�}U��z5sy������z��w���� Z�X�N�{��P�����U�܏S������xI�����j�=� �C@4���o�6E��ԷR917���l�5���v�*3��_S5�t'+=?�$��wB8�#��8��9]�y*�5��{f�	״�i�r�i�%S�rà�,/���������֬C�D`]����f�aZ��2�Nښ.��'#���
��D��jH��xd+���O�VA�����T��1�����K����=�I�QA��ɕ�Ϸ�'%X��u��g���c�paz����I�[�����^�Y�X��w�'ؙ���pKɫ�^�h�7����?^$���1��������%X@C�ġ���q\-�y�[RLVR��y�a�\�Kh1�%��D7����]7���8���5-��@8/r�^���hX%+M	ĵ��ͮ5�)[8sZ|�k��%���7[z~��Ja�ʱ��x֏×sh�K��yb�;�# �����@��e2%��hA�`�9U�t3���$�еH�=�/o�͔
���c�.f�	�nVl����м��WU<$N,5��	5H����8\� �uA!D�93�j��]���?R:21/���;�{���5jz��G�����#�澻|��u�SEK�(�ev��!F�%b��4c�ڵ0��t/S���:8���T%1V{*~P��Β��KFΜ�#�E�9�w��������[R�M�汶v��J4���oI�Xi� �r�N����cNUrԡ�)�{B~4�@p�߅%�ާ+�Ҭ�n�k/�h;�v���~2�)�����*	��[s��1�$��[�<g�c��ʮ���(��o�G:��<�Gr�TDq����ޒ���Lq\u�^���7��96�)�����u\)(�'�G.y������i��|�Ժ'K���y�"`C�5	��bD��d{W��ƌ�,r3Ź�>ʙ�E�u��ŗf�D�ٖ��i����r�W���J	POT���l��� S�H�G9UN5��#Rѥ�N�A�ǃ���A� �T#��UHCP'=3�}�R_�b�7�T��V$ؠ֝���J�5���nA���[N�2�����I�D`�.��ߊ��"����3c�F�)�o�ٸ��c�)�#�$�%nwn��峝~:�@	˾��h&I����"�1;w�f�"q������G�{�6���5f�?0 찪�e�Km���i�sl�VYڊ�V0O�ē�9 =Y�j>�{=�MZ��s`-���b�@�4��ӹqR�	l����A�.�\�Ԧ1��ͻ=YM::5'�$R�w�t���  ZI��	�cR�1/�AQ� �"����.N]�-`��Z��ދо�I{P�;��3�2���:�,-	��3��5�vt�K�7
�CN��e.�jݾ�'��yYtt5BԎTPKwf�����<���$Yl]�_�Y~�#���)]t��"�[QP�-W�V�y��J F��(8�ۨ|Js�1���ڹ��")�Faz�7yM�S��&�ߋ��2��2jR��D,Z
��/���zT���/
�B7�W�1ُ8?6�-��a6���+�fOdl�%��DSoq6��g�"ǹ���}`�oQt2r&�qPqP?�I�~c?TnI��x����j�7�	-Ծ���2�L_��5�����b�[��1y�l#H�`�&R��������_[V4�ɷ9�WS2�:��<(����)�Ns-��Ė���,�2"Y�)	����H��5̤�Is�!��xH���×�s�4Y�+*�4��P<؀�W�bw����ʐn�W���| o��Ф�gS��o�Y����[�G����>B�[�K�ZE]���\���ǯ�)GG���ɨ�#�r��u,���s��0\��Q����+�8�y�^��n$�ґ��XiRj�܇���
� so����e��B^�E�>:{�B�i�Y�-^�7�H�����\��%�$к�[����{�[�X;�#.�/k������ji����
	�I�$E���l�?b��9E����湖�HA�K��9���Q���*bu�cZiU�o�D.���[�Z�z=*e��Ey�QG��LA�Gh9�}G+z�ǋA�&5��O�5�O�X��=�v
��?��´s��5~�Vԣm�_��DA�?���H�A>_.I���@��ƏNR��@Un#��ha:!���HFYn)I}�RZ��Zt�{uS�����M3�{I8�NB��A�f,��[�������5�z����S|(�l���!��꣊ųE48�{ez�ҫ�N�����1&�l��vpx��U<W[�#支 ��:5<5�ޤ{����eA�h?���Y��{}mp��Bp(�O1Vd-k �͐��8oտO\�P���Թ�F�M�4�g�h���78�����!++�z1xL؆��$P_eD�O�w�Tl%%�����¼ƒ�j�4wV[�Ӑ�X�c+i<FGb�߈���/�Z��=�|ֆ��|*N�SU.�W��dE7sc3��mf��ʌ��WCQψ	��$���TI�6ElI���h=O�!�����?�b'�̴�����ӡ4�������땄j�~�s����g���dD�.l�em��}����'�"ʹO���m��أk��U���^�����I���J��!� CV\,��#��su���!��E|V��4l�v���_|\���wU��Ɔ�.a����C@�:��>�4c�J��;9_�YԳ�AfBԎ��i�Y"��˴+|�]��ݪz����L)H-���^�^Kup����[�DSrL{C��()l��'������:�;۞ٻ�������� 1�m���dj�kw��8��1��q�����<{���H�Ǿ$�'�I0!�������m4�)[���T�Mj���py�d�)	D��#�	ē���$F�8>��({ B��RN���q$Ό����
y��p)S���`�n�؇�̠�l�J{��	�_�'�dʣ�޻��S���]XbG���;8z����j
�H���5}�o]x�e�'j,Ʉ�H��>�͊\$OC�������ꭚ�6�wRCm/�$�̃Ia������ڦȯxJBø��N?nqD�1���)��Xݽ���YH���w�R���˦�ƪnz�9��gK�p�#�y�36%DZ���+" ;���S�@�]a6K`��E������CnY�AY�2������-W�L`Lk`μ��m~�6ZB3Tĳ�wI{S�m�ǈa�]�&���h���޵ ��;�U��B'�  �<�+r�Y�ġ����+�)G1��=c��&@@w���={����v�#'�S��~4��iD�7Q��s�����j�8�F���O�֩l|�M����ڰ;i�����<VptR{�V�������SLr4&�����;�kޖ}�J�c;S�s�h����)j��N���/.i�7��>b�"�=�s��h~��wo����d]�]�YYwV;�X�F�q���jf	x-���޲��	��X$b�� ~w��bHH>��C�\j���M$�PΛT[_8p�J���'J	�,���'���Yz陎���&��R4d�_�G���z�;M�3\��ÉZ���OF^��q�d�������xSQ���Ũ8J�,�B隣���z���z����zE�/�D}p��9Yr�I�`Ӹ
�IYR�؁ @#��z�1�\��x`�R�:�p��F~!��n�'��!�}��R��?/d��;z`��"j�`l	.Z<8����
H)��t3�w�]3���}CN���������l��(����jn�%�>���B��7�ڝ�6��!�����ϫ�IB�����RA	�����L��CY��k��s����A�&��"����l�#���(�^e�Y~1ԏ���W85c��#F���>GU<�ғ�jA����'�1&�-s-�뽏���̔ɇ$"��9��4���4��^��IE� ��n�U�؀'h���'Ը�J��J?9�`f��qjf�-��!��1\ZqA�v)a�'�+�n�>No��ަ:`2�9�]�JA~��%f[��S(��*%���^,�O���oE�R�>Wة�߭��d�4>:���K�bT�9%Î�dh��d ���mbj>��m�w�Y��+���rAg4x9J����S/Y!N�{y����"5���-{�ө��5��@ w�%�P�߁�+u�0��k��lT��v��] ��m+� �)�o��z�!)}��_��͵���pc9�gUNQ���t�<h� W��rĐ�&�$���B�����t&jHL��&��m1@���M�)��5���zB��4�n.5k5Y�	����?֟x{1�y�?&��}~���v��z�p��.����|��ފX��%%�S\J�O������z��͉�R@��cs���$a���Ԕ�"c:�Q�1�΍寔5;��n�ո����!Ve�n��bSc����N3w3���xQ���Rç��Ic�*�(ʢJ�����4uU�A�S���K�S�����vɳ��<���s�Mu�=��Q����x�{��v�He�̣�B�Ӌ����\ Y�x�(��=��}��g�F��:/1ƆO���ΞW�|E��$`�
sح��^y�R�[A�'�D��ʃ�!6�Q�Dr��ԐAYD0��ǜ>��}���*(�a��%�b�����S5	�=F��qrC�fo�.�6��ZYC	�*KH�����d�3��<s��Sb7�n��ʽ��S�2%r�ؙ�����sB��_ތ,XD:��R�KbZ9!~�����VT�R�q����U?ⷾ��K���;���K7SP��n�ut_(:���e�/�'��+��R��JՖ���}���K% �kn$<�C�T!�����Fj�9UQw���r�I�4]�x9���� �U���~��x��k��������MrR��?��^#�e�?EP�D���ܮyr�E�ak0�4ےS<$��_�������KzE-��_e��
@�MQl�ˈQ�"'6M��� [��(�	��փ�Tgq|�nf"��2������{��3��mo�TtS!�fI���c�I�b)[8{4��Ӡ��ھO'�HE�Bx��:�3�I���%l����f�u�} 	YsW���h��%�yb�ݨ���M�{���r�U3	s��t��)�x���ޘf��r̰s|K9�H���C3l6-m^I�O�-8&��f�ӵz�ޕY��{�{�`K
�˺��m�M<�+m�1+���u^��E�=(���������m�dr���~����t�DzZDh_Z��~����pE�u�?R�o��&L^��:��;-(�4S�ߋ���!����~W�b�)�4�؊����Clᨔ��w�<�V��n���@|�;�*��ǈzCh���ni���a�%'^s{�&+�L����\�}=`u�f��8 �6�k_-�2A���0�bMw��l4����:�ߕ�QMO�"���b�s\��+K^]ɫ��,	k�6㚊�i���e"�XZ�2Fю?��9���XU|���F 6�VA��K�G�^]�6�O-B18*sE�K��?�aNR;�AF���\i��ٚ`�ܺ��qb�T��������Tԇ����6֕��]�A�z�#�+r��#�u@$q�������ư�w(q��K�aQi��|�S�A��t��d�.�G��+h����)r㈇�6 �*.��zsO~����*�nE��xx�lt���c�l�W��PǠ����,�}o؀^���-+aaj��:�L]M��7�s3��!�~��ˎ���?���(`>��n��B[z[�#RFU��tvj���낹Y�jA.`sw]����� � ��������%����"=<��9[w�+��6[�W��փ�4Q	�L�1�V�,tRy���
|6�H\ߘ�OyR@C3�'����뽒!i�=�x���vcE0�plp�Æ�P
k7'����4Jb���:Ex������B�)b7 �R�Q�Q���k=��O�8#����a]�TM+� ���Ib��U��*]�.v��Y��nN�8d�
������E�t���K��)3G�[|6s�8�d�x�F�!EM��"���S-?rm�o��k��x�O%'�k��3Հ;��XĹ����p���v3tRI@/�u��ƲwxĬ
��A�����`I4%�K�.�н8_�	L����K�zm�Q�ޒ�R��7�;�2��k�� ^0~��o���4�"�2^B�T���[1"��
�����#۳,b!�#��S�m�˪�c6�U�Z�.�]�&}�%&�.;2�B¥��R#X�,W�-Jz��8��-�� ���܎z�}������҂Ky�/�:�5B>����9��$k�5C�����J�}�o���Z�x���+�T��i&q�.k\��1���4��c]�hwC.̻P��%�vo�q�B�!c���~�� &��>��