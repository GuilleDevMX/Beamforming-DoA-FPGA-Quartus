��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V���T6�I!b�����JL�9E:xۯ�4C6���`4�P}���	%�BT�o�s~��3�qr�{�܀��V�yP�!UWw��^��ʧj(�����	%�3_�9_�S�FJHW��cpG��<䖺���~�PCI�6�����g�3@z4�y�JY�R2���lF�@�Ϭv�b1{k���!M���ί���5�8��"A�QPp����YZ�@�|��R-��A��bx'�cLϵ`"m�
�A�> Yn��j֨:C\|�GJj`R�)���p������B`�R��>LX7�K(+ۙi'�!���h��dî���W��q)`A�!��;6����7�	6i�L-�5��T�}Ŷ�m�)�س�k�Z��U쯶��s�9-p-��$�{*۴��@BMm�&!\c��9/���J[�¥�{$�)�YKB]:�N���\�/b�	���[��bt�ܸzO�cWn�L>�؆�!�ԸrO���AD��S��`t*	�;p��X��Q��W����~4�9���D�n!P�u�,��K�}kV1thz�>��(�E�g|W\�>e�K�#x��p��ĽE���~��`�-��/ ��WNJĆ� �n<�8x�O~�5}�>�(#�`��B=w�Zǉ0���_B��(�'�8kE�CbY�Q���JD�8_��pT�(�B��+(?�@Q�gh'ڻ�%������ŬC�Q����I�+��-	��FQ��V��*R5�h*b8<]B���-7�� .�Q�J΅hru%�Wu�H�)�q�H�cx{��g�3�3�c�[�d���^�Ou&��X00���6iL�^�]�B�HÌ�tS��
M+�6��s�4Ө�̃���L��45�w�A\m���j��H�>��7˱�9�(r��U1�Q9�3F����]�W�k�<$�Y�����' ��OУ \�|
�?�%
�H���d%RTp�uA$<z��_y3��K�BA�.g�Sİ��_(.ܝ�ɇYS��4��1hdR���3�-I{�b�ɢ}Jj�لhm�1d���hG�m�s����P��؅{�cwl2i��n�rq�P��FL/�a��B6�����w���#�}h�\�K� v-!_��h�7��`Wlu���բD�]� �p��VU;��/�Xh�<v���V��xN�SM-q�s�1�^_8Ƶ�N��g�l�s���У��&&�s��VR���h������u�h�(��;1�_0冄y����Ths�@)}�-mw�b���	*ҡ�]{

����;��{�ҏ}�!���e�S{��
~���$��W���+yg�×ƥ���j�4��8&�T|W�	@0��dU�K���@��X���;�O����S,A̚�T�$%r��������
B<q�9"�Fx�#o�½�7`��@�'鹛2�"�!#�<T4K62W�M����I;�lA!?�V�C�褝�x�o���IE]O����3B�p�0�����x���;c��E�J������聅��6�UY����\�>����x�6�ɺZ��.�*<3Ŧ���1�;��#m��
4�遌8��ǂq��D��8�ۢ��<�ހ1�jL��X�����ȃ�k> �tB��o>`��Qp���T�ҧ.��?u��CѤ�/�Ҏbj����%z��9@�]+��O&l�I>^^U%ݿ���h7$;�8�iZ�[g�p��U|��9Z%���H�m��
��,���4o�Ȑ]��C��~�UC�P�W�Q ���q��-��� �������:�������ӆ9C:�lf����n�3=�˼%�Ǎ^��i�L�-��e�3�~�T�.�����Y�����r`���ٕ���|���49i)׍}@�d��2)lW�)�;;���s����[�E)�>�&�(���Rd�S��}*%/��cc�[��{u��r���
D��e�QG��[�ۃ����}�&�<E�����Ǆ����<�����_��8����(�
� F������;�^�i��l��tN04�G�Q.�Gp��h��3��)�T�����9|�ʆ~%����E^�� �ӖB����94혓"!�Є����r,��S2ѱ�.u�c�Y5�6�Q*��|�C�乙!�8�C�I_�Bc*>/?�=�*fu����D�V$�guӤ��l9���`x�E{6��	�{77g�t�0\�9���a��*�6��p��5~��;բL��6�G�բ��O�Q�*�r�����.dU���B:��D���� &�L��7���]x}�����0+���L�#h�6��b�&���(��-�l-TвP4x�t�+J*KL�����YN�B����v�ý��VT+�B�ɜ�b�"亶�VuMHZ_	.7�o!ο��fY�(=��r0��1�F��.K�%0T
��]裩jO8K�*���{Ir�{ϑ^󨕦Ҧ��~�x;e��T*��>?�:붙�׭1�no�`
�=�w���(?,�#����)<?�9f�����q��MP�o7��f(=�貄�DP�Y��{�F��A����$3x.13J��xt1�M{"Zeq�=h
2�����2~g��R֗�(���|��{;�6�	�?���Ɖj|��&[�Y�+"HH3�B�!2�tf��{|�r��:�җ���j�(�/.�S�m����~�� �;��e���N�A�.�?�bP�(���+D���P�u�Y	0�a��]���х8%��rЁ�zg/�W��x�t�,K�_8*V@ʻU�0�ް���_�C�����1��0=G�<Ol:K��p_�O�[ ��!@7�k��9q�.o()���::��`XL�0���p�G&
��$"/���~������)�M�,��2��+�� P�!U�\��[lu%���{���-}Z��3�:S:�S'���M�� ����=��E��t��#=���y�=K�
�@j�fb��9iy�m��Fwi���)�x�ǧ�d)h)^�L��}.l���x|lw����P�7�n�#Q���y%��Q`�*�BWyΖ޺��yJz[�r��J}�flވ�S�ռ�|�|�i/����]K�mH�9�xr����,q�F�ͩ����k���B|�5�$ʢ�Q����S ��Y����S:���Y�/]ҧ���T�ra#�WG%�L%����~�*���ƶ悔d	e8���]�UU�'�F��q��+I��3�q��=��w���CJ�Gm� m�0�dB���E���<Peס;�P� � Dr�k��@��&�����0�wK��$ſ�sW��\�4}|�
-	?Ip ~� �櫭�r_�l����Bۇ��+n&�Xd��I
L�$�m,�/Ip�QK�8&(�a*�cr���tj~���S��R��"��u=��ߵi�2��O����ʘ�T��}m���$gT�VR��t#Ԩ��ˑJ_w�����k_鴟�
��ΙҤC�@�~�&��ċxFW��Dpk �aV�'>_q���}<�e�]p�C�M
 Yl^9]0Q8�8Up����٧���)v����]�bo��N�����D����)W�:�42V�]L���/��Z�醤D�4�hI$.f
w���W}�!&��֒Ee���׵U���[��IUcۥf�ʈX?����7\]�uQɨ? %�~�ɋV�- ������H����K�ڸ��Eز�}<;��?��I�񝐺�,�t�V~��	E�I��6&��OO���YNǘ!$ o�֌%]�l��d��!Hq/�t��zJ�k��H|=L�)о�b�:�)���-�_����)|�*�N(2�A��.�%`m���^�7���L�O ���4k[�����>�&��0&-�,ōJ@�׶i�z�r�::�g�M��ͅ!��B�O"����O}�L?�qj���P��jP%��$wz@3�J3����EY����L�N���e����c��[�0ɜʒ�����>���\'�����,eŎ�GNoamN Y�ʈ�
|���� ���2
�V���"�Dȑ�� ���DC�beҙc�Mt�p�Ţ��M���+J{|%­��}M_�����\tr�d�Dr2-�;������D��ዒ���Zw���:a�Ov@y���l�'�|���س���:��z�#h{�֨�#��|!��H�:e}[����w(QE?�n���ǻ��a��"cW}�"ĵ��N,U[M�j�Y*����z�}�� �Fb����i���ve��63���/N͛��?��w�p+�XZ������֢��>�`��PU���E�[O��C�s²R��F�.���Ћ