��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���~�`���sB�U	Ù���iCK������F~��y`�N��D��wx~�Nz�#d��(/#�V��:�t>74���ϥ<W�e�a*b���.}U0������L�)����M�V�-lq�P�b<��Ө������Y���#���Y|z<��s��lb�� �8|�=L�8y�u"���lT����Ni �`&a@l�?����|�ַ3{-�*ٟ��(�>|�=?�n�ܴ��=\Sޝ^Ҟ�%�`ߴ�d����q2ս�r��D�k���Wa#$�Pq;���I�y��h���>B��;�m�rt��I~��mJ̦���0���Bdg�9�	�����V)qd@&�D��$�f�1v�1��$*1�)u�����N�)�b\U����� I�?c(h��0�Wh��O��-� /�{{	�y�ڡ���X���ɞ������1�����öv��Of�:̗]̮�����6j�8�4�����[�{����S�L�ߓ�!��r3��n
�0F�0PSr�&;�L��3�s�g���]���rWY�c�������:#�����l����>X��`è� �����[v7��b���}�g�yv�#Ԩ���f��E@n�	?Y�� 1lD�5m�qNg�gκ��2�9��V�VTL�1�S�b�\�����'�AG>��[(]x��zi3;V�[{<0��]�n����y�<Q�6�>;�6��	���%n'=��jrK�:��UpF`<�M�sLٽ�����=������r;��Q��9����EXh��$ώ�� ;��M��e	}��_Դ�^��8���s������}&QNG:�j*r�i S.���m2��k�'��M�!G�æ�i�<ج���l�YLߓ�$rL�.b�ܱ�= pn��i����h��2Eh��zo@~afijJ���c8aaEf�r#������t�j��lk��.�!�J-���%�fY�g?*5ʢ���*�������T�Ҽ�A�Z/F��ǔ��_yz��@ID�1S�*FgB��C�j�P��e�K撘	#���}������.y��rxH�Q䗛�~�$5A�A��c��0���cj'�L��
dN1×߯�ߞ$c��v��$ ��gQ�O��|������V�������ԡ9 "}���J�������	ˣ̕[�Uc�啍����Q'�
.�3����4��>�x�|��}�<����<��P_�`)L�R�:y�-����_������}�Aez�Q\� \rG��C)4��������杳�K���H����a�M,��^M�_���WFN-��BSGn$�����*^y�k�BS�0)�#č����@����Z�l�OP����LN(K@��@��x�>�{�@��K�}jJS1�|����&����0��P\�kvU@zǶ�Jf�&L�'$H$&]w�ch��ك����i�죸*��7�f��[^��4,QehN�M��B�d�� ��fs��O7�sh��@*l����ET��T8��7��_� �!<�2§�}�[#B\�F� p�/E�Ne�u�=l��3m3,ȉ��Y0�������?L���3`#,�B���h�R6$k��P!���{%��$��*�d  VC�kPi1�8�w���� �/�����f̤��!O�;(Q�N
J�[T�VK��t���Ʈ���u��Nd&����q�1���� S
�`�̆���y[m�[��0)o��n�$f�|����=�!ɫ���t�</]�*���Ɠ����3L�J�``÷|���LR����7:� ����nŴ,�ܴ�S샱\A ө��Nf`��I)\%��������n�w����'�Rrxv�O]���v��<V�j�ȚΟTOmN�h���x>WBF6p9sfWH��1}���<�/�VE	D>W��}��(�=uK��j~\��L���dS����e���)F7s��h���FϚQ�f������T�L>�1�|�p��Aυ㫆�|�:ٖ���6ɼ� �I�c���H��=�rcf��1�6j�]��=	���\�h!�� 	A.�ai�;��d� �u�	���#ナ*��