��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈڽ�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��*1��x��H�8�����ʴ�kX�CY0 �Ɖ�����r�|�g���-�"�lköi�-�V�;��uc�p������(�?ք<�������v�tI/i���`�l��K� `���i�	��^rf���������(�r�[�3Y�Դ��#��a����"3�Ty=Ҫʎ���cG�������~��|��]�1�?��X�
���?J�\z���(���ëٹ����"#�3������RG/1���v>�vu�+��� 	�u*�ǩ�0Շ,�=@��Q�t`��ϵ�5�N�pi�#!�u������d
�ҵ��W��	��.Jd�
o7D�	%+�xUƓH�q�,-�_��|p����	(%=���v1�_�����@~D��������B��)jT����$ἓ�"�����&�d�;m�[(�?���گ��/�^M��`Z���xP���	�%��-D�hb]��`9���n��������ϩpe����z�k�q��>(�����|��<����1������M۰C1���EJ�����1V� Ii�x�),�T����e�����F�%z��!�����5u�#�3��m��"?�r�~�ƮPX�9�w2dM%�cX�}�2Յ�ԩ��$��9�0 9A�
K����BO��5� �e+L�-sN*���ώ�T�^��f�=��a��]:����J���3��pBC�
+t|��ϓ/�,�����Y���>c8b>L����Z�~���Q�k	%�������,桺'�� G$.��R`.�ùh�Lh�N�A��.@���nU$Wnj@wC�����ڥ�`�L�E2�� ���{.3D�B�]8�[���1��6DS�6��mk=8�#��8c�^R@�fvj��af�SMo�"�$���;3+,R����ģ��p6�촒��E�ֽ��L��q#���>�d��4���y���������FU��ǚ�����Cuֵ�恩]�}�����b_'�{9�u��� D	j}`Q�H�!����?�E�c�d o��^�٢�t�^0p�ی������Z0DL����#���qץ���'���}���0�H����x/5����N��I�j'HڻyK ~]��g-*)K�ϗ�ò6z���?�E��
����m`�<�֦d�AF��J�� �d���'�r��?8�y���b�F��qd��@ޝ��!�v��Z��@�P�^[�i��������s�y|5��'oʰ��V���H<���hR�L
+0���X�Pl͙3N��it��FQ(�X��)��E
c�5]�x	�FAo��&�#5������1��;~��:�����f�e3����v� �Z�����0m����/����i���'�w;�4���ZIf��o�R���ה����8{��g߹DlG�۝aޠ�7!/�I �a���5[�r%x[8�t�D[Y(��V��,9.�s��J�|��h�"����Y�4{s�r���X'��N�F΋]љ�����7��z��+�Hw��p� ��w����t����#d_�啣�?P�g�ϼ�7�- �7�˹;���0�cHK	�5p#�y���E����������QB�=DG��������1��r��;�`h?v�	"{��1 Gc�$L�[0��Nd�"�u�������=C�Ej��k<ϛV���X[j���FP��0UH-mLX���q|P�Ws'���va�b�����N3���h�$���j�j�����{=�L��O�Q�B���J� �0;9���B����VL����_cr٫�������7q:�Ci%�K��r���Ӂ-�:,16J��r�zSn��c;���e�n�}���bcX�g��K���l>N`G�<Ǣ��B��*~�}�z���c�~,��Rh1#*f�p��+��R���'_
m^S�y�~������KS5,�@��P�?��[Q�bD� ����>s	�qeU�v�m�P��Y7Ԏ�EC���6��Ӆ������"Ǐ܄�zK+OE�v�׌V��QDu%�J���u=�תQ&#b)�lJ;%��Gw+j�/$<i�$��F�uO�8u�V�|��zĎV�S$��'x�'�_Xpu>�Xl�rh?�St���'�Io�nƺ��S0�a�3H��f�t�I?k��?w�5�B��
������n>5h�;ޜ�Cb�
ܼ��}���&��ӭ}�\"x����8^-�7�� �hi� 0�W��Ƹ���*79u����ۧ��)v�(�3��fC�8�Ꝙ͍TN#�QmS���ïD��QG|k΀#�x� D^��ZU!;<��ۃ>��&ȢPU��Ȍ�SF��٣N�f��'@/��j�\�}�4���=.�Ƈmv�L�]�M�z)*�� ,|[7�p��"�Zm��ͮ�+�C���^�Z�6b�A�����L�'��ݰ�*�3����NMK�ʵ���=�%/L�+��H)���r�[�Y��ga�r�q*�]5��@�܀��':���S
� "�5��u��%+L�ie�H`L��Nģ��s�yG~	v�0U����XE*[�'�>W)�&�8
A��S�{�4z�P�-p�Li@m����� 0���j+���M�D3�!'>�r�Jx� ��k{w'��8r_#�E]�u9�x��L��'���!y��mg�[2F��rܭ|��قGC�>� ������:�i�p�w\������.�B?�7�ш����������;p~���@��l�2��i�'�&��@;�nJe^z(��$�F<��pP����� ��bTAP(�n�:B"#�݉�ӄ�������B'LD�z�\����I*6vV�u>� w�+B�O(W��n���n���vEn���Y���RPf��m�@�α���w��Tb=�,HCR��$o8t�r��Z��������a�$�>����א'����4!,֕t��[�ΐ�0��Q�����⋛I�?gn7�2�n�
�F�Oo�-��&�L�
���r�:%};�3��(L�0�W&�u�Sunx���xyz}x��� ��h�m�<0ӹ�h#�F�7݂˂��=�R�![�
>�zm�F&�Q�K��Ԇ� e�@f�g,[��3�6&2�(��+��+�w1��=
���e[GS�x�U�i|V�s��v��+��˲��
K"q�X'B��7)?^��>TbFWy��il����������#���8�W����I�Zօ�q�%QF�s�<��n�e��KiW`�n��0�y�6���ؚ�{�&�$�T0?�-�U3Kx�nxjڑd,�?�)����J�?�~��߉J��76���}h)�W�Wr:-�����d���涱K)5��S��~m:v��wUu����0��J��Cd!1�{QEfd�z^�m�cg��C<�:�Z���#ӄ�~Y?�OG�w��x{2������&�HQ�7��uv�չ=)7���I��P�sư����`\��6�,�" �\�[N`H�*5��X#̶���-�-�7��sE�]k�CЂ��墉���u���k��pH�4%�~N�V�3�k+3�zZŉAX��l����g�YL��U�`��u�qX�	/O��:��p��b�\J����e �#��p�U���'3:P���D
�u��2ˌTE�D���j�4��O�A7%9�[�"MjTޒ��	��JP�Ex�ZK.��rN��,g=�Gm�(������ 1;�Ӑ6�!�����4tiH��=*��S��r˅@T0�gNW�:�=��*m��\�_ �+���q_�iM��3��s�F��ʧ4�r�;���t<�O� ��eI�1W�嚄Z�%x����k�Y`�-"�<j7��a-�%����l�cW�����a�؀ϟ-��i\��LO~�e.\�(�<{�o[oW��6�It���W��!��##�b^�ZO�#�5����Y��g���D��M�	@�ꒄEN����m��Z��n�tX���o~ؠ�����u�£��%t���6=��kX��d���g�z�-�PdM.�8a�e7����4���*�d�PN�:7�P��DC����;��qB����(
LU�{^��L�CK3�D�{|�1��y%�f�oI�[�F�����R�Q�K�k��Us���G���K���|r�M����0����y�P+=*?�(K7L�q?}n��D���f'��.�u���4��hr�ָ��	�y���%��sn��ډ���<n��V�[�]L#<W���O����c����47á�P�Ͳ_Ǫ��
��3��B�'�b���k��� ��L&���yOx)`����G��jh��`����Bij��w��&�ς`Ur�Hc�?���;M]�t�
���1<��H����u��`�aT1�o+�����S{䷂!*`��c��"�(��P�#���U���y?`�'^	�M�Rf4 H�5�#п;�{ڤ62���qM���4�v�R���{�+��#�#sc>�Q��z4䔤G(�<��񣊝-�mɟ���=a:^
��_I)���a�qE6p��WVMx���K�m����Q��h6Rw;��-ZB�dx�C�fGߜ���&�z�[)�u���!�)��ݐ���4�R����?G�Ғ4�f�E����*�v�S[p�X��LA,�QOK��!I��}RKw�sU��5��ӴW����ók�:���Lͻ�-Kh]�b�EV�����遉Fy�D<.O��K� &�2���d��8��'~�=�z�]�0r8�gRI��� Z��p��C����Mٖ�W�o��O���~�?;�E��G�Y�@�y����!`��
��_�۹��Ӈ��&c����V"���ǡ
&�o���,����Ő�6���"��=���B~Yam���vBp5�_��_`!׋c��{F��<+�&c5<4�!q��x0ۏ���=�g���[A���{e*a�w� �s��%�� ������mc�{�VQ�N1��YX���LO����7�LX����?�����B.�E��i<��,�r���W��Ꙧ��HL���w'{���S�hoX�7�=���H6�F2��EN�@�Ʃ�X��IK[L�0����'� 
^K���gbP����<��L�@���7�4�y��:�����Cm�O}�N�v���WK��]Zы���rJ �<�6�b����Y�UO�l(+��q�y؀ޭ$��u�3�=��?0����OeNt��W<A�n��/��I �*%¶�s�
Q�4�:5"Y?A3���T�*z��za!���nz��W�x�*�o� ������ݴUiCz���Z�� *c?.`'��Y�	��V&�'�$��Z��ď\�\�b6I��IL=�k�s\ |����P_��?��m�w��ҭ��y�a�kp>ݫ>�e�xbp�=�ߴ���G�.�u�_e6��Z�B�g��˒b��eG\H=�r�P����<����#�G�a�A{,�]4�g/p�ngp��#D�̓O�z	v:_�s��{�y�Gg\�i�����;�U��>^I��6~�(�[�=��L�I��6����A6=>ԟ��J~F���=q:�2��[��٧)ږ !r'��\��c0�V5�����%�Vo8Y}}1��<�N4E�ow^�E��Y��ʉ®��8MX;��\��@�"��~ݹjw�dc�,�i8ClU���p9��x$Њ�O���e����TÛGLz�?	��"�dW����	Ҙ�����ݴ�	M7�hT�=��AO��:�����aFĀ�����hB�7��{'���`����D�1�d���g�W6ɱ���F#ASo��r�Rl-W����h%�F6�����`�/#nG��v)?�I]xzr�$���*�!GA���B@Ҏ�9�J �����B��� w�Z�x�^'|���8 e�@ս(Ad��t'`�XL��ײ�C{�[��q�)�:���Dl8�m�m���~���>�/C��� ����)�S��!����8����T��-�i�qe1�m����j�E1�`��ZrW�ܺ�pjQ���*�+� �ꮦݛ��
D�aY�f�z������z���*tRyd*)L��*
���=sjZUayǁ���-�o��[0����7��Y �q��<���h�ѹv0uQF���#S�W����#ߧ����a��t�{;|,�6� �vs֖	#��Y���(�
�y���^�Ͼ��]�*-���l�92���A���L^�!�`��c�`�%������j��y8�厪����ķ�v�+�}�}���\^�+��V�2jc�'�{u��*��èn���L:��'���a��ha%�����E�����)e�9��{k��k����������J�K{I�C����>���a���;Uu��<�-.�����H�iQj��ĥ�o������G�;�:pmBSZ�OC���p<1=�}>�hX�h4&���7��jBPN
@�������k����[�������[��ov V�L�b�}Hg��Αq�cmP�j-(�*�M������!c�RMtn]��Vִ,���f=P�jX�Q����Z���ɂM�!�;����F
�k�_{I8����8v���: p�!�^��9�.��oGB[(o����̺n25D�Q�_��o��*�c3c��⺹�~��a�qYm,��k��oW�+�<?�;�*�Up�I2ŕ�5�[R���p��*��ܯ�~W	]���97��������1��Xl��@��$��LMD��>D=0��_�>k����$
��]J���������ꡛj���CF�,��a��|c�6��[�cT��:F؏$�=7Yfu@�������
`�c��$+"��������ѩV�%��}st�Lu�4Gs5P�� >��Du{���RI���7`��N��K�����X����e�n���Sv�:F�S)�)�G갎�B�F	zp(�8.L�)� 4d�=/�/}?���x��ǽ}L]Q���ag,C�N~�wY�u�\��p12���6@8�2k�S�ȷG�xE�|Uف݂��5,�ׅ�H��?��,9��!��0ݾ��+RM��>�B�Y�2��[r�ܷS���VP�ا{��cx��{�p�d���!Wy-�(mu�q'
�.�t(� L�,R��G�R��F뎎d�-�'+�6�w��!'����9�(f���u�O���! ��'Sx�q�Dl��(�ϛH[����'���n�'�rv�؋e�dvM8�縿����GT�c��l1�Y/�K��D�I�<��㝛?&���sϙp$�`o[n)mȆ�k�q�0��:��n'6i@��h|QN ao;:����'e�{��w<l�;K��D��?(A�R���u�G�6_����C!_�ss�-�"v�d�:���"�PXQ&����(������Rf@U"k��&���~��یP$�m���wR�қd1Qb�T.��+�Lȭ��6F-	�3����f�����Q����|X,�Jh�MK�_Ö����;��?�l$�@��U9��7å�0��A}�B�5
���2>ܟ2&O��.H�P�n��������5��D�Z�t� ��2ec�DT<�4����R
���۞��a)B���$��e���<�l��R��1©�AZ���O)
9����%Qe�B�qN�}�J%1���S�@�	(g?I�n��X�,d�T��
��8��G�"
�Q8��DN�l�dQgL���,��)�$4��/ZbR�,���Cay�����I)���h�譬�~��_ϒ 挢�>�<�.hl0\�U`q�v$�L���y*��X��*%-L/���\l�_#Ydit�+O��Y����*��,%��H#�a�R2��'Q�8{��P~�h��A�q�F�?֭�p��[��I��d��1�sE4��f�� a(y"�� ����6j��	�`b����Z���ᐳ4DAEŚM;|ʙ�z���@y��du��R���؆=�Q����$=��&�1�J���=���P��]-����j���N}/��ݲk����������a�ҩ3���Unf��e�U�#!Ml^g��iV�"u��s�3E:�E_��k���V����;{�ޯy�~獅����t1K!�DL]7��?V����<ʵo�^�e�2�tC��}K�����:��l	/����%.D��a(8f�D��ͽx�A�����5�,����i�H�9G+|�Y������
b$1)R��=.�jM&7T�3xT���ܟ�k�	�E�+UF�Y�ćJ�����Z�W1n�e���q���"���T�	4�y8���q��&���W�+��,��3箮+߉<��p�C�_3<�8�鐔M
y�� W���E���[y�l`jR0��.R�[�H�c�Y��9�c�g���g�қ�%�&�W�ikk��R�u���<�Fv��,�)�+�e�׆��)1kl��t�*�Kj]_W��-��ʂ8�4��v�O%VU�ͧM�03�G�S&q�����k�@�R\�V>��;�50g�Y�/_����÷
��8���>eNX�{ͺ�V�,����^���=�f��Ԥ�p�uRO����G�zVz5��c*��&I�u��SœOKK[^[R��B��AT�T)�x`�ΕpG�BM$�M0�K9XK��3��{`m�ր�I����ʆ�ށ0T/��{�W������s�!��6�}o�����/�e˟oD�P���m��,s��y�Y�Ŏ�n"�Z��Y��؇Ҳ>Q?o�fE��
��s�Ni�Ě�7���)�N���3Guj;���,��qq7D�y�2�ow�%�3�C�-��K)�"���TN��*.���0�Ր@���(
�%���&���ז�f�:�TWb�J�y�Lk�<	��m*ݯ>�GT�PvWK�|� >�&t���R�1��Mnc�x�A�-{Ӭ��CF��rac�<�w�gC�Gy�y���:l�������(S��.�5�Qc	n٬��ye5OA�|�|��rQ�/����x2�w�&�@�o��X�G��f��]܆�����.j�����ل��E���*x?G�^�O&�3�ޢ���i��JI:7����Xb�D��ƒ�bDk���H2?�f|���UH�V�6H����9�Idi�S�𐽆K5��y�9���V
�s6�F�޿\i����/R�� �sw�{Z��)�|'O�?S��=�XE���wz�\�4�xd�$mR�1��w�d]&N[��Fn"��<�o%j1|��X���:Xc���Xѽ�Fo��Q�������;U�d#�t�qjZ��$��/ܮxh��2��&��)hPM�?3�p�8JBW��+�K�����Y�������3`�����Q-)�$�T��M.
q��bE��� {.ˑ�FC�nkS��(��m�zբWv<��ND,:h��o�*�����Bٍm����ƀ7���w�\�w��)��'k�W���i;�uf����D���<�;��,�2��ht�A�%J�oT9t���	פ�	aVd|_�/�}�#���j]�!+T-�<VQ��rJ���m�H:
@ppl0"��v��g���c��gK6��~����0"ٿ��h��`y*.�O'�����-�$��L�Zr�<��(bH�N��ŝ���a��jp1��]@�%��Q�^�)˩o&�o���y���}O/��2�5%���>b'V��v$�Rc��C�{��t��o�4�D���ǃE�H�C���dщ�����=�,ㄳ���!@B �^s�
�;)��=�A����
H $�[����Sjdo�,\�~���9fA�!{�U��]�{�!=����a�*�4[nbm�
;��rR� AMT��V��a������WH%�\v���2t�O��<h��7��Ep��(2����2R�ާ� ���ې�����q=/�>���!���)a��x�14G#�x�/��?�JG*�VM�fP�ɖv�7��q7��E�������	�zA3�����İ��I7E� �<ŊG	��E0e��qa���aO�|`���9�E��`�q���u"r�Fc��nkٸ�R�Q���	^�A��ш>c�%��m��dG�(��Y�T��@q"j_���i�Nm|��H���r�C��Y �+/B��>��������a)MĀ�Dt0�c��j�f%���Ù��1_���8UW=L*�u�V�;��g�_q�C��H�F��i��y5"t\3m<�ę�<B)��2M0��Wn��_ Ot߭]�qo����{����z���5�s]��Y5�+��]��<�Ι��.���[9��Z�~�r7ȷ�Im���;���R6é�tK����5��7��^�������H�E	ir�l^���9>`p>�!YI6��W!�S��s�f�f|��N<���׎h8 R�q��26y�lg�I�����i�{l	c?�}D�LԴN�+�_e�*J��`pLᳯ_/n����D�X�}�l8�f�ȏO�)�{��I��:���GECŵ��/1@���/88�[/�|hl�r̰�y�C)��5(<���W��ڵ�i���#�j������%[�#,���T<9��0rt���w�ۊc8?`�����?%!Ү�F{�D��!�ʻA=��򼠒[ �/[�"���5�n�����``������Yi߱`�S	r7�π��s���Y[��-6aۇ�߷b���{��\��\dF��*kZY��p�V����+�1w�Y'QM�]`|����Mxһ��:ψ�Ť4�I&��DvQ}��O�cy�@���?��G�#�c(�=��/�-�͛���,�N����toǅi�������@�'$�K?G��@��kqk�͉�-��j=H1��D�h2��]�C	V
℠ô�r{d�g�U*ZX�m�֑�4'F�J�Qe/��*f�?z�N�eSQ_��v�z�1H����B���
�w��x�
q�2��%���!����՘�6��/��=9��гi8�Nx���l��Ȓ�f[����4���|�h����	�з��I��[�b�q��<�S��[���s�Gg�!@��<��E�^���Ҫ'�����&�Y��S��B�ƃ=��5�bW"$GfFJ�?v��ZGG���D���|G��3��rw�W�{IE�� ���Z��?���K�_r�����S/OyIC�" �O�u���,��І��|�?�N�0*RA��[Zz�z($~'�����ъ��^�М�4v%�[�ˢg�&�z" ��m��洼��>��֘�w���nh��:�I�K1�X������te�2KZN�6VӾ�v�?��P8��V>��>ؓ I���#<һx�%�Nh�F�Y!��V2��;?��a��j��xjؿ;eg�����.ݔgЦy�3,��3a�#/����px�ߤN��t��#�"��My}���[(gʜ�b��#'��g�Rg�8(��AX�dj?���L��|Ŀ�!�U$����U�5���*�|r�����Z���+H�"k��5͂p��m|�0�k9����66۲W��L`E��
0w�hU�ݬ�a�B����`'�`�
2��8�#�CY��둻�?wEX/Hx3r����۠m�FՆx1��W{��J�k��I:��Wd o�|��J�Fʪ�~����� �>P���&o6�%?���1��c��*SL$�5t���������}��	���1�j"jv<���G�J��in/�xZ��?M��=��5������Z�J��*�� g\�BZ�_��A�/�%�.VB��]d��}v$Vs��]ٯ��T7��ډ�_�������-��nPS��&��-��η�^Q[g�A~/�ڨs=g�t�HI�{�q��!ފ���O��Z󴁖;HH)�\�}��nyZ4���vm�������%*�L�ǯ�b���=� ��v1V'AO�C#���|��OƏ��W��w��A�I
暱�n�@�@ͳ�j�L��5���G�(�`#>C�r��CkZ �`M�2����]�񊥈�ܲC�Gߖn��O����7�Z�^R���ڧˢ�l�o���2�I�XY�$�2���W}v8[�,NZL5W"t̍�E����!M��3�ػ�¥�L���ޜ����A�cK�/at.ᘬ�a@�E������ m��A�F��Y)���[W���ጕ/8|���������C��)>x�\t�c(�KJj��qV���1r0��D�ǘr<�u2��%w�@���i�S��/!%[�K��E��B�u�(�����R�eAwYt��������b'�j�c.k��)��D�)蟷2�Q4.p��X�V%w��p���Ih��?@b�ҟ;�?�ڴ`�׾�I�w�jS��� -ُ0������RO�-�����F���7|����]�r����c-V/A�Hs>���e ���@�w"���v|�u��⩖JY�a�>�e��յc����d�u�a��[�M_�*�v�
��y��(��:Y����