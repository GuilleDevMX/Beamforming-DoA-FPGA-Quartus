��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��z�ٖ��"�a�Nc�	QB[�.UK�̿�t:��-!m���9-:�@�.0��U��譌�^��R�}/r��� |sQX��6��?�kˡ��!WXq?ӈ�-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#��U3�q�p��*S�^�b1T�m�A9��V�������$�[hɄ�gl�(5��1ˍ�R�)�]��w��k0�cʮՃ,^4��#�S�/,q=�U>��+G�N�!�k�7&h�![�/
8Ĥ ���cϡ��*�~�rx�p8;.��]�Ǫ�{B���ʬ�������2����Ԑl���7��~Va�憉P��e4MВ?!�4gᆹ*Y�[D���M;��r�L|��E_0��Kc��כ��w�_P�G<�P��&c @��P	�u.Y���:��2�Pd���E�>���%�1BfݹF�9�W��
�Aa�d��Q�YԳ`H�&>sUT�GM��g������r@R�|Gd'ie�=p��3fJ4*G��[ƃ1���OA���u3�r����:�k,��av��c��`S-���3L�!R����q�Ul�7���h*H��eN����(:����]]�r(�/�ހ��U_~�=� }��z�g��*ڟkZ.Y�y�)�-+��R<�����}���|&q���_�[>��[��c_t��TW8�I�[>[�ov@mT"ك��kaej�h�]j��ѽ����D�]������+��Lw��o:l�^Xi]l�Ƈ�����z�:��O�f'
�O�s�<�˲�]����XuN�T�q('��pG9����,+ڜH����N�,yQTP�w��&����e�*�)�_ɱ��.�ЙQͫ�:5���Fq�r�ڐ4���'�=fM���I_�@r��;.��Gb���c_��J(�Wl��Z������:��1QA]���"�}��ګ�ۏ�Ե`ӝZ�3A���M{S��u_�����l�����y6��~����3�\0�֘�_��=�E*c���d�\p�,���p�t��c���Dv�UwY0c�W�X���?��TЦn�]�S��j�TE�Ck���ױx5K�6�=��f�n�@1�.~�ZX�I�Ҟ����.��CW�\�A�Ȅ�Yx�BE�f#���ۯ�[!��@��9���9[|3Ofx~���&�F ��?��`���O�]��Fè�ƭ8a���p&��2A=�9o��(ܨ�F� J�@m���"Ci�Y��O8?��u�6��q�4�cy,g0*@w��=�k0b���ۘU��߯^��8=UTZy��kY��21P>��Vղ���л�r�L�\K������������'��A��p\u{Jb��lW
0��$�g�X���4�teI�{����ǯv"���Ŕ�3i�s�Kd4�d�����#Zt�~�(t��&��u}
ڥU�#!�����n�D���)�A��d�G̬��!�2�ó^kJש��AKi�U
���1���:����x�8	O"rú�H[�4깅�{ݥ<�`��0	g�d�p���J�}��\Kx7~C�_^��fk��ICA�|Gk�hȩ ��ip�L��0d�O^�f2X&����d)��糨��r����Ї��$=f7Ⱦ������,�